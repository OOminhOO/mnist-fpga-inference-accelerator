`timescale 1ns / 1ps

module tb_cnn_core_top_time;

    // ========================================================================
    // 1. ��ȣ �� ���� ����
    // ========================================================================
    reg           clk;
    reg           rst_n;
    reg  [7:0]    data_in;
    reg           data_valid;
    wire [3:0]    decision;
    wire          out_valid;

    // Loop �� �ε����� ����
    integer i;
    integer err_cnt;
    integer c1_cnt;
    integer p1_cnt;
    integer c2_cnt;
    integer p2_cnt;
    integer fc_cnt;

    // �� Latency ������ ���� (�߰���)
    time start_time;
    time end_time;
    time latency_ns;
    integer latency_cycles;

    // ========================================================================
    // 2. DUT (Device Under Test) �ν��Ͻ�
    // ========================================================================
    cnn_core_top u_dut (
        .clk        (clk),
        .rst_n      (rst_n),
        .data_in    (data_in),
        .data_valid (data_valid),
        .decision   (decision),
        .out_valid  (out_valid)
    );

    // ========================================================================
    // 3. Golden Data �޸� (Hex ���� �ε��)
    // ========================================================================
    reg [7:0]  mem_img   [0:783];             // Input: 28x28
    reg [7:0]  mem_conv1 [0:1727];            // Conv1: 24x24x3
    reg [7:0]  mem_pool1 [0:431];             // Pool1: 12x12x3
    reg [7:0]  mem_conv2 [0:191];             // Conv2: 8x8x3
    reg [7:0]  mem_pool2 [0:47];              // Pool2: 4x4x3
    reg [31:0] mem_fc    [0:9];               // FC: 10 logits (32bit)
    reg [31:0] mem_pred  [0:0];               // Final: 1 value

    // ========================================================================
    // 4. Ŭ�� ����
    // ========================================================================
    initial begin
        clk = 0;
//        forever #5 clk = ~clk; // 100MHz (10ns �ֱ�)
        forever #4 clk = ~clk; // 125MHz (8ns �ֱ�)
    end

    // ========================================================================
    // 5. ���� ������ (���� �ε� -> �Է� ���� -> ��� Ȯ��)
    // ========================================================================
    initial begin
        // ���� �ʱ�ȭ
        err_cnt = 0;
        c1_cnt  = 0;
        p1_cnt  = 0;
        c2_cnt  = 0;
        p2_cnt  = 0;
        fc_cnt  = 0;

        // (1) Golden Data �ε� (�����)
        $display("\n[TB] Loading Golden Vectors...");
        
        $readmemh("input_img.txt",  mem_img);
        $readmemh("conv1_out.txt",  mem_conv1);
        $readmemh("pool1_out.txt",  mem_pool1);
        $readmemh("conv2_out.txt",  mem_conv2);
        $readmemh("pool2_out.txt",  mem_pool2);
        $readmemh("fc_out.txt",     mem_fc);
        $readmemh("final_pred.txt", mem_pred);

        // (2) ����
        rst_n = 0;
        data_valid = 0;
        data_in = 0;
        #100;
        rst_n = 1;
        #100;

        // �� Latency ���� ���� ���� ���
        // data_valid�� ó�� High�� �Ǵ� �ٷ� �� ����
        @(posedge clk);
        start_time = $time;
        $display("[TB] Start Feeding Image at %0t ns", start_time);

        // (3) �̹��� ���� (28x28 = 784 cycles)
        for (i = 0; i < 784; i = i + 1) begin
            data_valid <= 1;
            data_in    <= mem_img[i];
            @(posedge clk); // 1Ŭ�� ���
        end
        // ������ ������ �ְ� ���� valid ����
        data_valid <= 0;
        data_in    <= 0;

        // (4) �Ϸ� ���
        fork
            begin
                wait(out_valid);
                // �� Latency ���� ���� ���� ���
                end_time = $time;
                latency_ns = end_time - start_time;
//                latency_cycles = latency_ns / 10; // 10ns �ֱ��̹Ƿ�
                latency_cycles = latency_ns / 8; // 8ns �ֱ��̹Ƿ�

                @(posedge clk);
                #100;
                $display("\n==================================================");
                if (err_cnt == 0) $display("   [SUCCESS] ALL CHECKS PASSED!");
                else              $display("   [FAIL] Total Errors: %0d", err_cnt);
                
                $display("--------------------------------------------------");
                $display("   [PERFORMANCE REPORT]");
                $display("   Start Time   : %0t ns", start_time);
                $display("   End Time     : %0t ns", end_time);
                $display("   Latency (ns) : %0d ns", latency_ns);
//                $display("   Latency (cyc): %0d cycles (at 100MHz)", latency_cycles);
                $display("   Latency (cyc): %0d cycles (at 125MHz)", latency_cycles);
                $display("==================================================");
                
                $finish;
            end
            begin
                #50000; 
                $display("\n[ERROR] Simulation Timeout! output_valid never asserted.");
                $finish;
            end
        join
    end


    // ========================================================================
    // 6. �ڵ� ���� ����� (Hierarchical Access ���)
    // ========================================================================

    // --- CHECK 1: Conv1 Output (u8x3) ---
    always @(posedge clk) begin
        if (u_dut.u_conv1.out_valid) begin
            // ä�� 0
            if (u_dut.u_conv1.out_1 !== mem_conv1[c1_cnt*3 + 0]) begin
                $display("[ERR] Conv1 Ch0 mismatch at idx %0d: EXP=%h, RTL=%h", 
                         c1_cnt, mem_conv1[c1_cnt*3 + 0], u_dut.u_conv1.out_1);
                err_cnt = err_cnt + 1;
            end
            // ä�� 1
            if (u_dut.u_conv1.out_2 !== mem_conv1[c1_cnt*3 + 1]) begin
                $display("[ERR] Conv1 Ch1 mismatch at idx %0d: EXP=%h, RTL=%h", 
                         c1_cnt, mem_conv1[c1_cnt*3 + 1], u_dut.u_conv1.out_2);
                err_cnt = err_cnt + 1;
            end
            // ä�� 2
            if (u_dut.u_conv1.out_3 !== mem_conv1[c1_cnt*3 + 2]) begin
                $display("[ERR] Conv1 Ch2 mismatch at idx %0d: EXP=%h, RTL=%h", 
                         c1_cnt, mem_conv1[c1_cnt*3 + 2], u_dut.u_conv1.out_3);
                err_cnt = err_cnt + 1;
            end
            c1_cnt = c1_cnt + 1;
        end
    end

    // --- CHECK 2: Pool1 Output (u8x3) ---
    always @(posedge clk) begin
        if (u_dut.u_pool1.out_valid) begin
            if (u_dut.u_pool1.out_1 !== mem_pool1[p1_cnt*3 + 0]) begin
                $display("[ERR] Pool1 Ch0 mismatch at idx %0d: EXP=%h, RTL=%h", p1_cnt, mem_pool1[p1_cnt*3 + 0], u_dut.u_pool1.out_1); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_pool1.out_2 !== mem_pool1[p1_cnt*3 + 1]) begin
                $display("[ERR] Pool1 Ch1 mismatch at idx %0d: EXP=%h, RTL=%h", p1_cnt, mem_pool1[p1_cnt*3 + 1], u_dut.u_pool1.out_2); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_pool1.out_3 !== mem_pool1[p1_cnt*3 + 2]) begin
                $display("[ERR] Pool1 Ch2 mismatch at idx %0d: EXP=%h, RTL=%h", p1_cnt, mem_pool1[p1_cnt*3 + 2], u_dut.u_pool1.out_3); 
                err_cnt = err_cnt + 1;
            end
            p1_cnt = p1_cnt + 1;
        end
    end

    // --- CHECK 3: Conv2 Output (u8x3) ---
    always @(posedge clk) begin
        if (u_dut.u_conv2.out_valid) begin
            if (u_dut.u_conv2.out_1 !== mem_conv2[c2_cnt*3 + 0]) begin
                $display("[ERR] Conv2 Ch0 mismatch at idx %0d: EXP=%h, RTL=%h", c2_cnt, mem_conv2[c2_cnt*3 + 0], u_dut.u_conv2.out_1); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_conv2.out_2 !== mem_conv2[c2_cnt*3 + 1]) begin
                $display("[ERR] Conv2 Ch1 mismatch at idx %0d: EXP=%h, RTL=%h", c2_cnt, mem_conv2[c2_cnt*3 + 1], u_dut.u_conv2.out_2); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_conv2.out_3 !== mem_conv2[c2_cnt*3 + 2]) begin
                $display("[ERR] Conv2 Ch2 mismatch at idx %0d: EXP=%h, RTL=%h", c2_cnt, mem_conv2[c2_cnt*3 + 2], u_dut.u_conv2.out_3); 
                err_cnt = err_cnt + 1;
            end
            c2_cnt = c2_cnt + 1;
        end
    end

    // --- CHECK 4: Pool2 Output (u8x3) ---
    always @(posedge clk) begin
        if (u_dut.u_pool2.out_valid) begin
            if (u_dut.u_pool2.out_1 !== mem_pool2[p2_cnt*3 + 0]) begin
                $display("[ERR] Pool2 Ch0 mismatch at idx %0d: EXP=%h, RTL=%h", p2_cnt, mem_pool2[p2_cnt*3 + 0], u_dut.u_pool2.out_1); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_pool2.out_2 !== mem_pool2[p2_cnt*3 + 1]) begin
                $display("[ERR] Pool2 Ch1 mismatch at idx %0d: EXP=%h, RTL=%h", p2_cnt, mem_pool2[p2_cnt*3 + 1], u_dut.u_pool2.out_2); 
                err_cnt = err_cnt + 1;
            end
            if (u_dut.u_pool2.out_3 !== mem_pool2[p2_cnt*3 + 2]) begin
                $display("[ERR] Pool2 Ch2 mismatch at idx %0d: EXP=%h, RTL=%h", p2_cnt, mem_pool2[p2_cnt*3 + 2], u_dut.u_pool2.out_3); 
                err_cnt = err_cnt + 1;
            end
            p2_cnt = p2_cnt + 1;
        end
    end

    // --- CHECK 5: FC Logits (Signed 32-bit) ---
    // FC ��� ��� ���� Ȯ��: u_fc.out_valid�� High�� �� out_logit ��
    always @(posedge clk) begin
        if (u_dut.u_fc.out_valid) begin
            // !== �����ڴ� Verilog������ ������ (x, z ���� ��)
            if (u_dut.u_fc.out_logit !== mem_fc[fc_cnt]) begin
                $display("[ERR] FC Logit mismatch at Class %0d: EXP=%h, RTL=%h", 
                         fc_cnt, mem_fc[fc_cnt], u_dut.u_fc.out_logit);
                err_cnt = err_cnt + 1;
            end
            fc_cnt = fc_cnt + 1;
        end
    end

    // --- CHECK 6: Final Decision ---
    always @(posedge clk) begin
        if (out_valid) begin
            if (decision !== mem_pred[0][3:0]) begin
                $display("[ERR] Final Prediction Mismatch! EXP=%d, RTL=%d", 
                         mem_pred[0], decision);
                err_cnt = err_cnt + 1;
            end else begin
                $display("[INFO] Final Prediction Match! Result = %d", decision);
            end
        end
    end

endmodule