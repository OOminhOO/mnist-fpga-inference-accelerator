module rom_16_images (
    input wire [3:0]  img_idx,   // ����ġ 4�� (0~15)
    input wire [9:0]  pixel_idx, // 0~783 �ȼ� ��ġ
    output reg [7:0]  data_out   // �ȼ� ��
);

    always @(*) begin
        case ({img_idx, pixel_idx})
            14'd202: data_out = 8'h54;
            14'd203: data_out = 8'hB9;
            14'd204: data_out = 8'h9F;
            14'd205: data_out = 8'h97;
            14'd206: data_out = 8'h3C;
            14'd207: data_out = 8'h24;
            14'd230: data_out = 8'hDE;
            14'd231: data_out = 8'hFE;
            14'd232: data_out = 8'hFE;
            14'd233: data_out = 8'hFE;
            14'd234: data_out = 8'hFE;
            14'd235: data_out = 8'hF1;
            14'd236: data_out = 8'hC6;
            14'd237: data_out = 8'hC6;
            14'd238: data_out = 8'hC6;
            14'd239: data_out = 8'hC6;
            14'd240: data_out = 8'hC6;
            14'd241: data_out = 8'hC6;
            14'd242: data_out = 8'hC6;
            14'd243: data_out = 8'hC6;
            14'd244: data_out = 8'hAA;
            14'd245: data_out = 8'h34;
            14'd258: data_out = 8'h43;
            14'd259: data_out = 8'h72;
            14'd260: data_out = 8'h48;
            14'd261: data_out = 8'h72;
            14'd262: data_out = 8'hA3;
            14'd263: data_out = 8'hE3;
            14'd264: data_out = 8'hFE;
            14'd265: data_out = 8'hE1;
            14'd266: data_out = 8'hFE;
            14'd267: data_out = 8'hFE;
            14'd268: data_out = 8'hFE;
            14'd269: data_out = 8'hFA;
            14'd270: data_out = 8'hE5;
            14'd271: data_out = 8'hFE;
            14'd272: data_out = 8'hFE;
            14'd273: data_out = 8'h8C;
            14'd291: data_out = 8'h11;
            14'd292: data_out = 8'h42;
            14'd293: data_out = 8'h0E;
            14'd294: data_out = 8'h43;
            14'd295: data_out = 8'h43;
            14'd296: data_out = 8'h43;
            14'd297: data_out = 8'h3B;
            14'd298: data_out = 8'h15;
            14'd299: data_out = 8'hEC;
            14'd300: data_out = 8'hFE;
            14'd301: data_out = 8'h6A;
            14'd326: data_out = 8'h53;
            14'd327: data_out = 8'hFD;
            14'd328: data_out = 8'hD1;
            14'd329: data_out = 8'h12;
            14'd353: data_out = 8'h16;
            14'd354: data_out = 8'hE9;
            14'd355: data_out = 8'hFF;
            14'd356: data_out = 8'h53;
            14'd381: data_out = 8'h81;
            14'd382: data_out = 8'hFE;
            14'd383: data_out = 8'hEE;
            14'd384: data_out = 8'h2C;
            14'd408: data_out = 8'h3B;
            14'd409: data_out = 8'hF9;
            14'd410: data_out = 8'hFE;
            14'd411: data_out = 8'h3E;
            14'd436: data_out = 8'h85;
            14'd437: data_out = 8'hFE;
            14'd438: data_out = 8'hBB;
            14'd464: data_out = 8'hCD;
            14'd465: data_out = 8'hF8;
            14'd466: data_out = 8'h3A;
            14'd491: data_out = 8'h7E;
            14'd492: data_out = 8'hFE;
            14'd493: data_out = 8'hB6;
            14'd518: data_out = 8'h4B;
            14'd519: data_out = 8'hFB;
            14'd520: data_out = 8'hF0;
            14'd521: data_out = 8'h39;
            14'd545: data_out = 8'h13;
            14'd546: data_out = 8'hDD;
            14'd547: data_out = 8'hFE;
            14'd548: data_out = 8'hA6;
            14'd573: data_out = 8'hCB;
            14'd574: data_out = 8'hFE;
            14'd575: data_out = 8'hDB;
            14'd576: data_out = 8'h23;
            14'd600: data_out = 8'h26;
            14'd601: data_out = 8'hFE;
            14'd602: data_out = 8'hFE;
            14'd603: data_out = 8'h4D;
            14'd627: data_out = 8'h1F;
            14'd628: data_out = 8'hE0;
            14'd629: data_out = 8'hFE;
            14'd630: data_out = 8'h73;
            14'd655: data_out = 8'h85;
            14'd656: data_out = 8'hFE;
            14'd657: data_out = 8'hFE;
            14'd658: data_out = 8'h34;
            14'd682: data_out = 8'h3D;
            14'd683: data_out = 8'hF2;
            14'd684: data_out = 8'hFE;
            14'd685: data_out = 8'hFE;
            14'd686: data_out = 8'h34;
            14'd710: data_out = 8'h79;
            14'd711: data_out = 8'hFE;
            14'd712: data_out = 8'hFE;
            14'd713: data_out = 8'hDB;
            14'd714: data_out = 8'h28;
            14'd738: data_out = 8'h79;
            14'd739: data_out = 8'hFE;
            14'd740: data_out = 8'hCF;
            14'd741: data_out = 8'h12;
            14'd1118: data_out = 8'h74;
            14'd1119: data_out = 8'h7D;
            14'd1120: data_out = 8'hAB;
            14'd1121: data_out = 8'hFF;
            14'd1122: data_out = 8'hFF;
            14'd1123: data_out = 8'h96;
            14'd1124: data_out = 8'h5D;
            14'd1145: data_out = 8'hA9;
            14'd1146: data_out = 8'hFD;
            14'd1147: data_out = 8'hFD;
            14'd1148: data_out = 8'hFD;
            14'd1149: data_out = 8'hFD;
            14'd1150: data_out = 8'hFD;
            14'd1151: data_out = 8'hFD;
            14'd1152: data_out = 8'hDA;
            14'd1153: data_out = 8'h1E;
            14'd1172: data_out = 8'hA9;
            14'd1173: data_out = 8'hFD;
            14'd1174: data_out = 8'hFD;
            14'd1175: data_out = 8'hFD;
            14'd1176: data_out = 8'hD5;
            14'd1177: data_out = 8'h8E;
            14'd1178: data_out = 8'hB0;
            14'd1179: data_out = 8'hFD;
            14'd1180: data_out = 8'hFD;
            14'd1181: data_out = 8'h7A;
            14'd1199: data_out = 8'h34;
            14'd1200: data_out = 8'hFA;
            14'd1201: data_out = 8'hFD;
            14'd1202: data_out = 8'hD2;
            14'd1203: data_out = 8'h20;
            14'd1204: data_out = 8'h0C;
            14'd1207: data_out = 8'hCE;
            14'd1208: data_out = 8'hFD;
            14'd1209: data_out = 8'h8C;
            14'd1227: data_out = 8'h4D;
            14'd1228: data_out = 8'hFB;
            14'd1229: data_out = 8'hD2;
            14'd1230: data_out = 8'h19;
            14'd1234: data_out = 8'h7A;
            14'd1235: data_out = 8'hF8;
            14'd1236: data_out = 8'hFD;
            14'd1237: data_out = 8'h41;
            14'd1256: data_out = 8'h1F;
            14'd1257: data_out = 8'h12;
            14'd1262: data_out = 8'hD1;
            14'd1263: data_out = 8'hFD;
            14'd1264: data_out = 8'hFD;
            14'd1265: data_out = 8'h41;
            14'd1289: data_out = 8'h75;
            14'd1290: data_out = 8'hF7;
            14'd1291: data_out = 8'hFD;
            14'd1292: data_out = 8'hC6;
            14'd1316: data_out = 8'h4C;
            14'd1317: data_out = 8'hF7;
            14'd1318: data_out = 8'hFD;
            14'd1319: data_out = 8'hE7;
            14'd1320: data_out = 8'h3F;
            14'd1344: data_out = 8'h80;
            14'd1345: data_out = 8'hFD;
            14'd1346: data_out = 8'hFD;
            14'd1347: data_out = 8'h90;
            14'd1371: data_out = 8'hB0;
            14'd1372: data_out = 8'hF6;
            14'd1373: data_out = 8'hFD;
            14'd1374: data_out = 8'h9F;
            14'd1375: data_out = 8'h0C;
            14'd1398: data_out = 8'h19;
            14'd1399: data_out = 8'hEA;
            14'd1400: data_out = 8'hFD;
            14'd1401: data_out = 8'hE9;
            14'd1402: data_out = 8'h23;
            14'd1426: data_out = 8'hC6;
            14'd1427: data_out = 8'hFD;
            14'd1428: data_out = 8'hFD;
            14'd1429: data_out = 8'h8D;
            14'd1453: data_out = 8'h4E;
            14'd1454: data_out = 8'hF8;
            14'd1455: data_out = 8'hFD;
            14'd1456: data_out = 8'hBD;
            14'd1457: data_out = 8'h0C;
            14'd1480: data_out = 8'h13;
            14'd1481: data_out = 8'hC8;
            14'd1482: data_out = 8'hFD;
            14'd1483: data_out = 8'hFD;
            14'd1484: data_out = 8'h8D;
            14'd1508: data_out = 8'h86;
            14'd1509: data_out = 8'hFD;
            14'd1510: data_out = 8'hFD;
            14'd1511: data_out = 8'hAD;
            14'd1512: data_out = 8'h0C;
            14'd1536: data_out = 8'hF8;
            14'd1537: data_out = 8'hFD;
            14'd1538: data_out = 8'hFD;
            14'd1539: data_out = 8'h19;
            14'd1564: data_out = 8'hF8;
            14'd1565: data_out = 8'hFD;
            14'd1566: data_out = 8'hFD;
            14'd1567: data_out = 8'h2B;
            14'd1568: data_out = 8'h14;
            14'd1569: data_out = 8'h14;
            14'd1570: data_out = 8'h14;
            14'd1571: data_out = 8'h14;
            14'd1575: data_out = 8'h14;
            14'd1576: data_out = 8'h14;
            14'd1577: data_out = 8'h25;
            14'd1578: data_out = 8'h96;
            14'd1579: data_out = 8'h96;
            14'd1580: data_out = 8'h96;
            14'd1581: data_out = 8'h93;
            14'd1592: data_out = 8'hF8;
            14'd1593: data_out = 8'hFD;
            14'd1594: data_out = 8'hFD;
            14'd1595: data_out = 8'hFD;
            14'd1596: data_out = 8'hFD;
            14'd1597: data_out = 8'hFD;
            14'd1598: data_out = 8'hFD;
            14'd1599: data_out = 8'hFD;
            14'd1600: data_out = 8'hA8;
            14'd1601: data_out = 8'h8F;
            14'd1602: data_out = 8'hA6;
            14'd1603: data_out = 8'hFD;
            14'd1604: data_out = 8'hFD;
            14'd1605: data_out = 8'hFD;
            14'd1606: data_out = 8'hFD;
            14'd1607: data_out = 8'hFD;
            14'd1608: data_out = 8'hFD;
            14'd1609: data_out = 8'hFD;
            14'd1610: data_out = 8'h7B;
            14'd1620: data_out = 8'hAE;
            14'd1621: data_out = 8'hFD;
            14'd1622: data_out = 8'hFD;
            14'd1623: data_out = 8'hFD;
            14'd1624: data_out = 8'hFD;
            14'd1625: data_out = 8'hFD;
            14'd1626: data_out = 8'hFD;
            14'd1627: data_out = 8'hFD;
            14'd1628: data_out = 8'hFD;
            14'd1629: data_out = 8'hFD;
            14'd1630: data_out = 8'hFD;
            14'd1631: data_out = 8'hFD;
            14'd1632: data_out = 8'hF9;
            14'd1633: data_out = 8'hF7;
            14'd1634: data_out = 8'hF7;
            14'd1635: data_out = 8'hA9;
            14'd1636: data_out = 8'h75;
            14'd1637: data_out = 8'h75;
            14'd1638: data_out = 8'h39;
            14'd1649: data_out = 8'h76;
            14'd1650: data_out = 8'h7B;
            14'd1651: data_out = 8'h7B;
            14'd1652: data_out = 8'h7B;
            14'd1653: data_out = 8'hA6;
            14'd1654: data_out = 8'hFD;
            14'd1655: data_out = 8'hFD;
            14'd1656: data_out = 8'hFD;
            14'd1657: data_out = 8'h9B;
            14'd1658: data_out = 8'h7B;
            14'd1659: data_out = 8'h7B;
            14'd1660: data_out = 8'h29;
            14'd2176: data_out = 8'h26;
            14'd2177: data_out = 8'hFE;
            14'd2178: data_out = 8'h6D;
            14'd2204: data_out = 8'h57;
            14'd2205: data_out = 8'hFC;
            14'd2206: data_out = 8'h52;
            14'd2232: data_out = 8'h87;
            14'd2233: data_out = 8'hF1;
            14'd2259: data_out = 8'h2D;
            14'd2260: data_out = 8'hF4;
            14'd2261: data_out = 8'h96;
            14'd2287: data_out = 8'h54;
            14'd2288: data_out = 8'hFE;
            14'd2289: data_out = 8'h3F;
            14'd2315: data_out = 8'hCA;
            14'd2316: data_out = 8'hDF;
            14'd2317: data_out = 8'h0B;
            14'd2342: data_out = 8'h20;
            14'd2343: data_out = 8'hFE;
            14'd2344: data_out = 8'hD8;
            14'd2370: data_out = 8'h5F;
            14'd2371: data_out = 8'hFE;
            14'd2372: data_out = 8'hC3;
            14'd2398: data_out = 8'h8C;
            14'd2399: data_out = 8'hFE;
            14'd2400: data_out = 8'h4D;
            14'd2425: data_out = 8'h39;
            14'd2426: data_out = 8'hED;
            14'd2427: data_out = 8'hCD;
            14'd2453: data_out = 8'h7C;
            14'd2454: data_out = 8'hFF;
            14'd2455: data_out = 8'hA5;
            14'd2481: data_out = 8'hAB;
            14'd2482: data_out = 8'hFE;
            14'd2483: data_out = 8'h51;
            14'd2508: data_out = 8'h18;
            14'd2509: data_out = 8'hE8;
            14'd2510: data_out = 8'hD7;
            14'd2536: data_out = 8'h78;
            14'd2537: data_out = 8'hFE;
            14'd2538: data_out = 8'h9F;
            14'd2564: data_out = 8'h97;
            14'd2565: data_out = 8'hFE;
            14'd2566: data_out = 8'h8E;
            14'd2592: data_out = 8'hE4;
            14'd2593: data_out = 8'hFE;
            14'd2594: data_out = 8'h42;
            14'd2619: data_out = 8'h3D;
            14'd2620: data_out = 8'hFB;
            14'd2621: data_out = 8'hFE;
            14'd2622: data_out = 8'h42;
            14'd2647: data_out = 8'h8D;
            14'd2648: data_out = 8'hFE;
            14'd2649: data_out = 8'hCD;
            14'd2675: data_out = 8'hD7;
            14'd2676: data_out = 8'hFE;
            14'd2677: data_out = 8'h79;
            14'd2703: data_out = 8'hC6;
            14'd2704: data_out = 8'hB0;
            14'd3196: data_out = 8'h0B;
            14'd3197: data_out = 8'h96;
            14'd3198: data_out = 8'hFD;
            14'd3199: data_out = 8'hCA;
            14'd3200: data_out = 8'h1F;
            14'd3224: data_out = 8'h25;
            14'd3225: data_out = 8'hFB;
            14'd3226: data_out = 8'hFB;
            14'd3227: data_out = 8'hFD;
            14'd3228: data_out = 8'h6B;
            14'd3251: data_out = 8'h15;
            14'd3252: data_out = 8'hC5;
            14'd3253: data_out = 8'hFB;
            14'd3254: data_out = 8'hFB;
            14'd3255: data_out = 8'hFD;
            14'd3256: data_out = 8'h6B;
            14'd3278: data_out = 8'h6E;
            14'd3279: data_out = 8'hBE;
            14'd3280: data_out = 8'hFB;
            14'd3281: data_out = 8'hFB;
            14'd3282: data_out = 8'hFB;
            14'd3283: data_out = 8'hFD;
            14'd3284: data_out = 8'hA9;
            14'd3285: data_out = 8'h6D;
            14'd3286: data_out = 8'h3E;
            14'd3306: data_out = 8'hFD;
            14'd3307: data_out = 8'hFB;
            14'd3308: data_out = 8'hFB;
            14'd3309: data_out = 8'hFB;
            14'd3310: data_out = 8'hFB;
            14'd3311: data_out = 8'hFD;
            14'd3312: data_out = 8'hFB;
            14'd3313: data_out = 8'hFB;
            14'd3314: data_out = 8'hDC;
            14'd3315: data_out = 8'h33;
            14'd3333: data_out = 8'hB6;
            14'd3334: data_out = 8'hFF;
            14'd3335: data_out = 8'hFD;
            14'd3336: data_out = 8'hFD;
            14'd3337: data_out = 8'hFD;
            14'd3338: data_out = 8'hFD;
            14'd3339: data_out = 8'hEA;
            14'd3340: data_out = 8'hDE;
            14'd3341: data_out = 8'hFD;
            14'd3342: data_out = 8'hFD;
            14'd3343: data_out = 8'hFD;
            14'd3360: data_out = 8'h3F;
            14'd3361: data_out = 8'hDD;
            14'd3362: data_out = 8'hFD;
            14'd3363: data_out = 8'hFB;
            14'd3364: data_out = 8'hFB;
            14'd3365: data_out = 8'hFB;
            14'd3366: data_out = 8'h93;
            14'd3367: data_out = 8'h4D;
            14'd3368: data_out = 8'h3E;
            14'd3369: data_out = 8'h80;
            14'd3370: data_out = 8'hFB;
            14'd3371: data_out = 8'hFB;
            14'd3372: data_out = 8'h69;
            14'd3387: data_out = 8'h20;
            14'd3388: data_out = 8'hE7;
            14'd3389: data_out = 8'hFB;
            14'd3390: data_out = 8'hFD;
            14'd3391: data_out = 8'hFB;
            14'd3392: data_out = 8'hDC;
            14'd3393: data_out = 8'h89;
            14'd3397: data_out = 8'h1F;
            14'd3398: data_out = 8'hE6;
            14'd3399: data_out = 8'hFB;
            14'd3400: data_out = 8'hF3;
            14'd3401: data_out = 8'h71;
            14'd3415: data_out = 8'h25;
            14'd3416: data_out = 8'hFB;
            14'd3417: data_out = 8'hFB;
            14'd3418: data_out = 8'hFD;
            14'd3419: data_out = 8'hBC;
            14'd3420: data_out = 8'h14;
            14'd3426: data_out = 8'h6D;
            14'd3427: data_out = 8'hFB;
            14'd3428: data_out = 8'hFD;
            14'd3429: data_out = 8'hFB;
            14'd3430: data_out = 8'h23;
            14'd3443: data_out = 8'h25;
            14'd3444: data_out = 8'hFB;
            14'd3445: data_out = 8'hFB;
            14'd3446: data_out = 8'hC9;
            14'd3447: data_out = 8'h1E;
            14'd3454: data_out = 8'h1F;
            14'd3455: data_out = 8'hC8;
            14'd3456: data_out = 8'hFD;
            14'd3457: data_out = 8'hFB;
            14'd3458: data_out = 8'h23;
            14'd3471: data_out = 8'h25;
            14'd3472: data_out = 8'hFD;
            14'd3473: data_out = 8'hFD;
            14'd3482: data_out = 8'h20;
            14'd3483: data_out = 8'hCA;
            14'd3484: data_out = 8'hFF;
            14'd3485: data_out = 8'hFD;
            14'd3486: data_out = 8'hA4;
            14'd3499: data_out = 8'h8C;
            14'd3500: data_out = 8'hFB;
            14'd3501: data_out = 8'hFB;
            14'd3510: data_out = 8'h6D;
            14'd3511: data_out = 8'hFB;
            14'd3512: data_out = 8'hFD;
            14'd3513: data_out = 8'hFB;
            14'd3514: data_out = 8'h23;
            14'd3527: data_out = 8'hD9;
            14'd3528: data_out = 8'hFB;
            14'd3529: data_out = 8'hFB;
            14'd3536: data_out = 8'h15;
            14'd3537: data_out = 8'h3F;
            14'd3538: data_out = 8'hE7;
            14'd3539: data_out = 8'hFB;
            14'd3540: data_out = 8'hFD;
            14'd3541: data_out = 8'hE6;
            14'd3542: data_out = 8'h1E;
            14'd3555: data_out = 8'hD9;
            14'd3556: data_out = 8'hFB;
            14'd3557: data_out = 8'hFB;
            14'd3564: data_out = 8'h90;
            14'd3565: data_out = 8'hFB;
            14'd3566: data_out = 8'hFB;
            14'd3567: data_out = 8'hFB;
            14'd3568: data_out = 8'hDD;
            14'd3569: data_out = 8'h3D;
            14'd3583: data_out = 8'hD9;
            14'd3584: data_out = 8'hFB;
            14'd3585: data_out = 8'hFB;
            14'd3591: data_out = 8'hB6;
            14'd3592: data_out = 8'hDD;
            14'd3593: data_out = 8'hFB;
            14'd3594: data_out = 8'hFB;
            14'd3595: data_out = 8'hFB;
            14'd3596: data_out = 8'hB4;
            14'd3611: data_out = 8'hDA;
            14'd3612: data_out = 8'hFD;
            14'd3613: data_out = 8'hFD;
            14'd3614: data_out = 8'h49;
            14'd3615: data_out = 8'h49;
            14'd3616: data_out = 8'hE4;
            14'd3617: data_out = 8'hFD;
            14'd3618: data_out = 8'hFD;
            14'd3619: data_out = 8'hFF;
            14'd3620: data_out = 8'hFD;
            14'd3621: data_out = 8'hFD;
            14'd3622: data_out = 8'hFD;
            14'd3623: data_out = 8'hFD;
            14'd3639: data_out = 8'h71;
            14'd3640: data_out = 8'hFB;
            14'd3641: data_out = 8'hFB;
            14'd3642: data_out = 8'hFD;
            14'd3643: data_out = 8'hFB;
            14'd3644: data_out = 8'hFB;
            14'd3645: data_out = 8'hFB;
            14'd3646: data_out = 8'hFB;
            14'd3647: data_out = 8'hFD;
            14'd3648: data_out = 8'hFB;
            14'd3649: data_out = 8'hFB;
            14'd3650: data_out = 8'hFB;
            14'd3651: data_out = 8'h93;
            14'd3667: data_out = 8'h1F;
            14'd3668: data_out = 8'hE6;
            14'd3669: data_out = 8'hFB;
            14'd3670: data_out = 8'hFD;
            14'd3671: data_out = 8'hFB;
            14'd3672: data_out = 8'hFB;
            14'd3673: data_out = 8'hFB;
            14'd3674: data_out = 8'hFB;
            14'd3675: data_out = 8'hFD;
            14'd3676: data_out = 8'hE6;
            14'd3677: data_out = 8'hBD;
            14'd3678: data_out = 8'h23;
            14'd3696: data_out = 8'h3E;
            14'd3697: data_out = 8'h8E;
            14'd3698: data_out = 8'hFD;
            14'd3699: data_out = 8'hFB;
            14'd3700: data_out = 8'hFB;
            14'd3701: data_out = 8'hFB;
            14'd3702: data_out = 8'hFB;
            14'd3703: data_out = 8'hFD;
            14'd3704: data_out = 8'h6B;
            14'd3726: data_out = 8'h48;
            14'd3727: data_out = 8'hAE;
            14'd3728: data_out = 8'hFB;
            14'd3729: data_out = 8'hAD;
            14'd3730: data_out = 8'h47;
            14'd3731: data_out = 8'h48;
            14'd3732: data_out = 8'h1E;
            14'd4246: data_out = 8'h32;
            14'd4247: data_out = 8'hE0;
            14'd4255: data_out = 8'h46;
            14'd4256: data_out = 8'h1D;
            14'd4274: data_out = 8'h79;
            14'd4275: data_out = 8'hE7;
            14'd4283: data_out = 8'h94;
            14'd4284: data_out = 8'hA8;
            14'd4302: data_out = 8'hC3;
            14'd4303: data_out = 8'hE7;
            14'd4311: data_out = 8'h60;
            14'd4312: data_out = 8'hD2;
            14'd4313: data_out = 8'h0B;
            14'd4329: data_out = 8'h45;
            14'd4330: data_out = 8'hFC;
            14'd4331: data_out = 8'h86;
            14'd4339: data_out = 8'h72;
            14'd4340: data_out = 8'hFC;
            14'd4341: data_out = 8'h15;
            14'd4356: data_out = 8'h2D;
            14'd4357: data_out = 8'hEC;
            14'd4358: data_out = 8'hD9;
            14'd4359: data_out = 8'h0C;
            14'd4367: data_out = 8'hC0;
            14'd4368: data_out = 8'hFC;
            14'd4369: data_out = 8'h15;
            14'd4384: data_out = 8'hA8;
            14'd4385: data_out = 8'hF7;
            14'd4386: data_out = 8'h35;
            14'd4394: data_out = 8'h12;
            14'd4395: data_out = 8'hFF;
            14'd4396: data_out = 8'hFD;
            14'd4397: data_out = 8'h15;
            14'd4411: data_out = 8'h54;
            14'd4412: data_out = 8'hF2;
            14'd4413: data_out = 8'hD3;
            14'd4422: data_out = 8'h8D;
            14'd4423: data_out = 8'hFD;
            14'd4424: data_out = 8'hBD;
            14'd4439: data_out = 8'hA9;
            14'd4440: data_out = 8'hFC;
            14'd4441: data_out = 8'h6A;
            14'd4449: data_out = 8'h20;
            14'd4450: data_out = 8'hE8;
            14'd4451: data_out = 8'hFA;
            14'd4452: data_out = 8'h42;
            14'd4466: data_out = 8'h0F;
            14'd4467: data_out = 8'hE1;
            14'd4468: data_out = 8'hFC;
            14'd4477: data_out = 8'h86;
            14'd4478: data_out = 8'hFC;
            14'd4479: data_out = 8'hD3;
            14'd4494: data_out = 8'h16;
            14'd4495: data_out = 8'hFC;
            14'd4496: data_out = 8'hA4;
            14'd4505: data_out = 8'hA9;
            14'd4506: data_out = 8'hFC;
            14'd4507: data_out = 8'hA7;
            14'd4523: data_out = 8'hCC;
            14'd4524: data_out = 8'hD1;
            14'd4525: data_out = 8'h12;
            14'd4532: data_out = 8'h16;
            14'd4533: data_out = 8'hFD;
            14'd4534: data_out = 8'hFD;
            14'd4535: data_out = 8'h6B;
            14'd4551: data_out = 8'hA9;
            14'd4552: data_out = 8'hFC;
            14'd4553: data_out = 8'hC7;
            14'd4554: data_out = 8'h55;
            14'd4555: data_out = 8'h55;
            14'd4556: data_out = 8'h55;
            14'd4557: data_out = 8'h55;
            14'd4558: data_out = 8'h81;
            14'd4559: data_out = 8'hA4;
            14'd4560: data_out = 8'hC3;
            14'd4561: data_out = 8'hFC;
            14'd4562: data_out = 8'hFC;
            14'd4563: data_out = 8'h6A;
            14'd4579: data_out = 8'h29;
            14'd4580: data_out = 8'hAA;
            14'd4581: data_out = 8'hF5;
            14'd4582: data_out = 8'hFC;
            14'd4583: data_out = 8'hFC;
            14'd4584: data_out = 8'hFC;
            14'd4585: data_out = 8'hFC;
            14'd4586: data_out = 8'hE8;
            14'd4587: data_out = 8'hE7;
            14'd4588: data_out = 8'hFB;
            14'd4589: data_out = 8'hFC;
            14'd4590: data_out = 8'hFC;
            14'd4609: data_out = 8'h31;
            14'd4610: data_out = 8'h54;
            14'd4611: data_out = 8'h54;
            14'd4612: data_out = 8'h54;
            14'd4613: data_out = 8'h54;
            14'd4616: data_out = 8'hA1;
            14'd4617: data_out = 8'hFC;
            14'd4618: data_out = 8'hFC;
            14'd4644: data_out = 8'h7F;
            14'd4645: data_out = 8'hFC;
            14'd4646: data_out = 8'hFC;
            14'd4647: data_out = 8'h2D;
            14'd4672: data_out = 8'h80;
            14'd4673: data_out = 8'hFD;
            14'd4674: data_out = 8'hFD;
            14'd4700: data_out = 8'h7F;
            14'd4701: data_out = 8'hFC;
            14'd4702: data_out = 8'hFC;
            14'd4728: data_out = 8'h87;
            14'd4729: data_out = 8'hFC;
            14'd4730: data_out = 8'hF4;
            14'd4756: data_out = 8'hE8;
            14'd4757: data_out = 8'hEC;
            14'd4758: data_out = 8'h6F;
            14'd4784: data_out = 8'hB3;
            14'd4785: data_out = 8'h42;
            14'd5276: data_out = 8'h4D;
            14'd5277: data_out = 8'hFE;
            14'd5278: data_out = 8'h6B;
            14'd5303: data_out = 8'h13;
            14'd5304: data_out = 8'hE3;
            14'd5305: data_out = 8'hFE;
            14'd5306: data_out = 8'hFE;
            14'd5331: data_out = 8'h51;
            14'd5332: data_out = 8'hFE;
            14'd5333: data_out = 8'hFE;
            14'd5334: data_out = 8'hA5;
            14'd5359: data_out = 8'hCB;
            14'd5360: data_out = 8'hFE;
            14'd5361: data_out = 8'hFE;
            14'd5362: data_out = 8'h49;
            14'd5386: data_out = 8'h35;
            14'd5387: data_out = 8'hFE;
            14'd5388: data_out = 8'hFE;
            14'd5389: data_out = 8'hFA;
            14'd5414: data_out = 8'h86;
            14'd5415: data_out = 8'hFE;
            14'd5416: data_out = 8'hFE;
            14'd5417: data_out = 8'hB4;
            14'd5442: data_out = 8'hC4;
            14'd5443: data_out = 8'hFE;
            14'd5444: data_out = 8'hF8;
            14'd5445: data_out = 8'h30;
            14'd5469: data_out = 8'h3A;
            14'd5470: data_out = 8'hFE;
            14'd5471: data_out = 8'hFE;
            14'd5472: data_out = 8'hED;
            14'd5497: data_out = 8'h6F;
            14'd5498: data_out = 8'hFE;
            14'd5499: data_out = 8'hFE;
            14'd5500: data_out = 8'h84;
            14'd5525: data_out = 8'hA3;
            14'd5526: data_out = 8'hFE;
            14'd5527: data_out = 8'hEE;
            14'd5528: data_out = 8'h1C;
            14'd5552: data_out = 8'h3C;
            14'd5553: data_out = 8'hFC;
            14'd5554: data_out = 8'hFE;
            14'd5555: data_out = 8'hDF;
            14'd5580: data_out = 8'h4F;
            14'd5581: data_out = 8'hFE;
            14'd5582: data_out = 8'hFE;
            14'd5583: data_out = 8'h9A;
            14'd5608: data_out = 8'hA3;
            14'd5609: data_out = 8'hFE;
            14'd5610: data_out = 8'hEE;
            14'd5611: data_out = 8'h35;
            14'd5635: data_out = 8'h1C;
            14'd5636: data_out = 8'hFC;
            14'd5637: data_out = 8'hFE;
            14'd5638: data_out = 8'hD2;
            14'd5663: data_out = 8'h56;
            14'd5664: data_out = 8'hFE;
            14'd5665: data_out = 8'hFE;
            14'd5666: data_out = 8'h83;
            14'd5691: data_out = 8'h69;
            14'd5692: data_out = 8'hFE;
            14'd5693: data_out = 8'hEA;
            14'd5694: data_out = 8'h14;
            14'd5719: data_out = 8'hAF;
            14'd5720: data_out = 8'hFE;
            14'd5721: data_out = 8'hCC;
            14'd5747: data_out = 8'hD3;
            14'd5748: data_out = 8'hFE;
            14'd5749: data_out = 8'hC4;
            14'd5775: data_out = 8'h9E;
            14'd5776: data_out = 8'hFE;
            14'd5777: data_out = 8'hA0;
            14'd5803: data_out = 8'h1A;
            14'd5804: data_out = 8'h9D;
            14'd5805: data_out = 8'h6B;
            14'd6293: data_out = 8'h16;
            14'd6294: data_out = 8'hC0;
            14'd6295: data_out = 8'h86;
            14'd6296: data_out = 8'h20;
            14'd6305: data_out = 8'h0F;
            14'd6306: data_out = 8'h4D;
            14'd6320: data_out = 8'h11;
            14'd6321: data_out = 8'hEB;
            14'd6322: data_out = 8'hFA;
            14'd6323: data_out = 8'hA9;
            14'd6332: data_out = 8'h0F;
            14'd6333: data_out = 8'hDC;
            14'd6334: data_out = 8'hF1;
            14'd6335: data_out = 8'h25;
            14'd6347: data_out = 8'h14;
            14'd6348: data_out = 8'hBD;
            14'd6349: data_out = 8'hFD;
            14'd6350: data_out = 8'h93;
            14'd6360: data_out = 8'h8B;
            14'd6361: data_out = 8'hFD;
            14'd6362: data_out = 8'h64;
            14'd6375: data_out = 8'h46;
            14'd6376: data_out = 8'hFD;
            14'd6377: data_out = 8'hFD;
            14'd6378: data_out = 8'h15;
            14'd6387: data_out = 8'h2B;
            14'd6388: data_out = 8'hFE;
            14'd6389: data_out = 8'hAD;
            14'd6390: data_out = 8'h0D;
            14'd6402: data_out = 8'h16;
            14'd6403: data_out = 8'h99;
            14'd6404: data_out = 8'hFD;
            14'd6405: data_out = 8'h60;
            14'd6414: data_out = 8'h2B;
            14'd6415: data_out = 8'hE7;
            14'd6416: data_out = 8'hFE;
            14'd6417: data_out = 8'h5C;
            14'd6430: data_out = 8'hA3;
            14'd6431: data_out = 8'hFF;
            14'd6432: data_out = 8'hCC;
            14'd6433: data_out = 8'h0B;
            14'd6442: data_out = 8'h68;
            14'd6443: data_out = 8'hFE;
            14'd6444: data_out = 8'h9E;
            14'd6458: data_out = 8'hA2;
            14'd6459: data_out = 8'hFD;
            14'd6460: data_out = 8'hB2;
            14'd6469: data_out = 8'h83;
            14'd6470: data_out = 8'hED;
            14'd6471: data_out = 8'hFD;
            14'd6486: data_out = 8'hA2;
            14'd6487: data_out = 8'hFD;
            14'd6488: data_out = 8'hFD;
            14'd6489: data_out = 8'hBF;
            14'd6490: data_out = 8'hAF;
            14'd6491: data_out = 8'h46;
            14'd6492: data_out = 8'h46;
            14'd6493: data_out = 8'h46;
            14'd6494: data_out = 8'h46;
            14'd6495: data_out = 8'h85;
            14'd6496: data_out = 8'hC5;
            14'd6497: data_out = 8'hFD;
            14'd6498: data_out = 8'hFD;
            14'd6499: data_out = 8'hA9;
            14'd6514: data_out = 8'h33;
            14'd6515: data_out = 8'hE4;
            14'd6516: data_out = 8'hFD;
            14'd6517: data_out = 8'hFD;
            14'd6518: data_out = 8'hFE;
            14'd6519: data_out = 8'hFD;
            14'd6520: data_out = 8'hFD;
            14'd6521: data_out = 8'hFD;
            14'd6522: data_out = 8'hFD;
            14'd6523: data_out = 8'hFE;
            14'd6524: data_out = 8'hFD;
            14'd6525: data_out = 8'hFD;
            14'd6526: data_out = 8'hDB;
            14'd6527: data_out = 8'h23;
            14'd6543: data_out = 8'h11;
            14'd6544: data_out = 8'h41;
            14'd6545: data_out = 8'h89;
            14'd6546: data_out = 8'hFE;
            14'd6547: data_out = 8'hE8;
            14'd6548: data_out = 8'h89;
            14'd6549: data_out = 8'h89;
            14'd6550: data_out = 8'h89;
            14'd6551: data_out = 8'h2C;
            14'd6552: data_out = 8'hFD;
            14'd6553: data_out = 8'hFD;
            14'd6554: data_out = 8'hA1;
            14'd6579: data_out = 8'h22;
            14'd6580: data_out = 8'hFE;
            14'd6581: data_out = 8'hCE;
            14'd6582: data_out = 8'h15;
            14'd6607: data_out = 8'hA0;
            14'd6608: data_out = 8'hFD;
            14'd6609: data_out = 8'h45;
            14'd6634: data_out = 8'h55;
            14'd6635: data_out = 8'hFE;
            14'd6636: data_out = 8'hF1;
            14'd6637: data_out = 8'h32;
            14'd6662: data_out = 8'h9E;
            14'd6663: data_out = 8'hFE;
            14'd6664: data_out = 8'hA5;
            14'd6690: data_out = 8'hE7;
            14'd6691: data_out = 8'hF4;
            14'd6692: data_out = 8'h32;
            14'd6717: data_out = 8'h68;
            14'd6718: data_out = 8'hFE;
            14'd6719: data_out = 8'hE8;
            14'd6745: data_out = 8'hD0;
            14'd6746: data_out = 8'hFD;
            14'd6747: data_out = 8'h9D;
            14'd6749: data_out = 8'h0D;
            14'd6750: data_out = 8'h1E;
            14'd6773: data_out = 8'hD0;
            14'd6774: data_out = 8'hFD;
            14'd6775: data_out = 8'h9A;
            14'd6776: data_out = 8'h5B;
            14'd6777: data_out = 8'hCC;
            14'd6778: data_out = 8'hA1;
            14'd6801: data_out = 8'hD0;
            14'd6802: data_out = 8'hFD;
            14'd6803: data_out = 8'hFE;
            14'd6804: data_out = 8'hFD;
            14'd6805: data_out = 8'h9A;
            14'd6806: data_out = 8'h1D;
            14'd6829: data_out = 8'h3D;
            14'd6830: data_out = 8'hBE;
            14'd6831: data_out = 8'h80;
            14'd6832: data_out = 8'h17;
            14'd7347: data_out = 8'h0E;
            14'd7348: data_out = 8'h95;
            14'd7349: data_out = 8'hC1;
            14'd7374: data_out = 8'h5B;
            14'd7375: data_out = 8'hE0;
            14'd7376: data_out = 8'hFD;
            14'd7377: data_out = 8'hFD;
            14'd7378: data_out = 8'h13;
            14'd7401: data_out = 8'h1C;
            14'd7402: data_out = 8'hEB;
            14'd7403: data_out = 8'hFE;
            14'd7404: data_out = 8'hFD;
            14'd7405: data_out = 8'hFD;
            14'd7406: data_out = 8'hA6;
            14'd7407: data_out = 8'h12;
            14'd7429: data_out = 8'h90;
            14'd7430: data_out = 8'hFD;
            14'd7431: data_out = 8'hFE;
            14'd7432: data_out = 8'hFD;
            14'd7433: data_out = 8'hFD;
            14'd7434: data_out = 8'hFD;
            14'd7435: data_out = 8'hEE;
            14'd7436: data_out = 8'h73;
            14'd7456: data_out = 8'h1F;
            14'd7457: data_out = 8'hF1;
            14'd7458: data_out = 8'hFD;
            14'd7459: data_out = 8'hD0;
            14'd7460: data_out = 8'hB9;
            14'd7461: data_out = 8'hFD;
            14'd7462: data_out = 8'hFD;
            14'd7463: data_out = 8'hFD;
            14'd7464: data_out = 8'hE7;
            14'd7465: data_out = 8'h18;
            14'd7484: data_out = 8'h4F;
            14'd7485: data_out = 8'hFE;
            14'd7486: data_out = 8'hC1;
            14'd7489: data_out = 8'h62;
            14'd7490: data_out = 8'hDB;
            14'd7491: data_out = 8'hFE;
            14'd7492: data_out = 8'hFF;
            14'd7493: data_out = 8'hC9;
            14'd7494: data_out = 8'h12;
            14'd7512: data_out = 8'h56;
            14'd7513: data_out = 8'hFD;
            14'd7514: data_out = 8'h50;
            14'd7518: data_out = 8'hB6;
            14'd7519: data_out = 8'hFD;
            14'd7520: data_out = 8'hFE;
            14'd7521: data_out = 8'hBF;
            14'd7522: data_out = 8'h0C;
            14'd7540: data_out = 8'hAF;
            14'd7541: data_out = 8'hFD;
            14'd7542: data_out = 8'h9B;
            14'd7546: data_out = 8'hEA;
            14'd7547: data_out = 8'hFD;
            14'd7548: data_out = 8'hFE;
            14'd7549: data_out = 8'h87;
            14'd7568: data_out = 8'h56;
            14'd7569: data_out = 8'hFD;
            14'd7570: data_out = 8'hD0;
            14'd7571: data_out = 8'h28;
            14'd7572: data_out = 8'h55;
            14'd7573: data_out = 8'hA6;
            14'd7574: data_out = 8'hFB;
            14'd7575: data_out = 8'hED;
            14'd7576: data_out = 8'hFE;
            14'd7577: data_out = 8'hEC;
            14'd7578: data_out = 8'h2A;
            14'd7596: data_out = 8'h12;
            14'd7597: data_out = 8'hEE;
            14'd7598: data_out = 8'hFD;
            14'd7599: data_out = 8'hFE;
            14'd7600: data_out = 8'hFD;
            14'd7601: data_out = 8'hFD;
            14'd7602: data_out = 8'hB9;
            14'd7603: data_out = 8'h24;
            14'd7604: data_out = 8'hD8;
            14'd7605: data_out = 8'hFD;
            14'd7606: data_out = 8'h98;
            14'd7625: data_out = 8'h44;
            14'd7626: data_out = 8'hF0;
            14'd7627: data_out = 8'hFF;
            14'd7628: data_out = 8'hFE;
            14'd7629: data_out = 8'h91;
            14'd7632: data_out = 8'h86;
            14'd7633: data_out = 8'hFE;
            14'd7634: data_out = 8'hDF;
            14'd7635: data_out = 8'h23;
            14'd7654: data_out = 8'h44;
            14'd7655: data_out = 8'h9E;
            14'd7656: data_out = 8'h8E;
            14'd7657: data_out = 8'h0C;
            14'd7661: data_out = 8'hAF;
            14'd7662: data_out = 8'hFD;
            14'd7663: data_out = 8'hA1;
            14'd7689: data_out = 8'h58;
            14'd7690: data_out = 8'hFD;
            14'd7691: data_out = 8'hE2;
            14'd7692: data_out = 8'h12;
            14'd7718: data_out = 8'hA6;
            14'd7719: data_out = 8'hFD;
            14'd7720: data_out = 8'h7E;
            14'd7746: data_out = 8'h30;
            14'd7747: data_out = 8'hF5;
            14'd7748: data_out = 8'hFD;
            14'd7749: data_out = 8'h26;
            14'd7775: data_out = 8'h73;
            14'd7776: data_out = 8'hFE;
            14'd7777: data_out = 8'hAC;
            14'd7803: data_out = 8'h15;
            14'd7804: data_out = 8'hDA;
            14'd7805: data_out = 8'hFE;
            14'd7806: data_out = 8'h2E;
            14'd7832: data_out = 8'h1E;
            14'd7833: data_out = 8'hFE;
            14'd7834: data_out = 8'hA5;
            14'd7861: data_out = 8'hBA;
            14'd7862: data_out = 8'hF4;
            14'd7863: data_out = 8'h2A;
            14'd7889: data_out = 8'h0E;
            14'd7890: data_out = 8'hDF;
            14'd7891: data_out = 8'h4E;
            14'd8321: data_out = 8'h11;
            14'd8322: data_out = 8'h2F;
            14'd8323: data_out = 8'h2F;
            14'd8324: data_out = 8'h2F;
            14'd8325: data_out = 8'h10;
            14'd8326: data_out = 8'h81;
            14'd8327: data_out = 8'h55;
            14'd8328: data_out = 8'h2F;
            14'd8347: data_out = 8'h4B;
            14'd8348: data_out = 8'h99;
            14'd8349: data_out = 8'hD9;
            14'd8350: data_out = 8'hFD;
            14'd8351: data_out = 8'hFD;
            14'd8352: data_out = 8'hFD;
            14'd8353: data_out = 8'hD7;
            14'd8354: data_out = 8'hF6;
            14'd8355: data_out = 8'hFD;
            14'd8356: data_out = 8'hFD;
            14'd8372: data_out = 8'h23;
            14'd8373: data_out = 8'h8E;
            14'd8374: data_out = 8'hF4;
            14'd8375: data_out = 8'hFC;
            14'd8376: data_out = 8'hFD;
            14'd8377: data_out = 8'hFD;
            14'd8378: data_out = 8'hFD;
            14'd8379: data_out = 8'hFD;
            14'd8380: data_out = 8'hFD;
            14'd8381: data_out = 8'hFD;
            14'd8382: data_out = 8'hFD;
            14'd8383: data_out = 8'hFD;
            14'd8384: data_out = 8'hFD;
            14'd8400: data_out = 8'h3F;
            14'd8401: data_out = 8'hFD;
            14'd8402: data_out = 8'hFD;
            14'd8403: data_out = 8'hFD;
            14'd8404: data_out = 8'hFD;
            14'd8405: data_out = 8'hFD;
            14'd8406: data_out = 8'hFD;
            14'd8407: data_out = 8'hFD;
            14'd8408: data_out = 8'hD5;
            14'd8409: data_out = 8'hAA;
            14'd8410: data_out = 8'hAA;
            14'd8411: data_out = 8'hAA;
            14'd8412: data_out = 8'hAA;
            14'd8424: data_out = 8'h14;
            14'd8425: data_out = 8'h84;
            14'd8426: data_out = 8'h48;
            14'd8428: data_out = 8'h39;
            14'd8429: data_out = 8'hEE;
            14'd8430: data_out = 8'hE3;
            14'd8431: data_out = 8'hEE;
            14'd8432: data_out = 8'hA8;
            14'd8433: data_out = 8'h7C;
            14'd8434: data_out = 8'h45;
            14'd8435: data_out = 8'h14;
            14'd8436: data_out = 8'h0B;
            14'd8451: data_out = 8'h0B;
            14'd8452: data_out = 8'hCE;
            14'd8453: data_out = 8'hFD;
            14'd8454: data_out = 8'h4E;
            14'd8457: data_out = 8'h20;
            14'd8459: data_out = 8'h1E;
            14'd8479: data_out = 8'hB1;
            14'd8480: data_out = 8'hFD;
            14'd8481: data_out = 8'h84;
            14'd8505: data_out = 8'h0C;
            14'd8506: data_out = 8'h85;
            14'd8507: data_out = 8'hFD;
            14'd8508: data_out = 8'hE9;
            14'd8509: data_out = 8'h0F;
            14'd8533: data_out = 8'h5C;
            14'd8534: data_out = 8'hFD;
            14'd8535: data_out = 8'hDF;
            14'd8536: data_out = 8'h1C;
            14'd8561: data_out = 8'h96;
            14'd8562: data_out = 8'hFD;
            14'd8563: data_out = 8'hAE;
            14'd8589: data_out = 8'hEA;
            14'd8590: data_out = 8'hFD;
            14'd8591: data_out = 8'hF6;
            14'd8592: data_out = 8'h7F;
            14'd8593: data_out = 8'h31;
            14'd8617: data_out = 8'hFF;
            14'd8618: data_out = 8'hFD;
            14'd8619: data_out = 8'hFD;
            14'd8620: data_out = 8'hFD;
            14'd8621: data_out = 8'hFB;
            14'd8622: data_out = 8'h93;
            14'd8623: data_out = 8'h5B;
            14'd8624: data_out = 8'h79;
            14'd8625: data_out = 8'h55;
            14'd8626: data_out = 8'h2A;
            14'd8627: data_out = 8'h2A;
            14'd8628: data_out = 8'h55;
            14'd8629: data_out = 8'h1C;
            14'd8645: data_out = 8'h8B;
            14'd8646: data_out = 8'hFD;
            14'd8647: data_out = 8'hFD;
            14'd8648: data_out = 8'hFD;
            14'd8649: data_out = 8'hFD;
            14'd8650: data_out = 8'hFD;
            14'd8651: data_out = 8'hFD;
            14'd8652: data_out = 8'hFD;
            14'd8653: data_out = 8'hFD;
            14'd8654: data_out = 8'hFD;
            14'd8655: data_out = 8'hFD;
            14'd8656: data_out = 8'hFD;
            14'd8657: data_out = 8'hE8;
            14'd8658: data_out = 8'hA8;
            14'd8674: data_out = 8'h35;
            14'd8675: data_out = 8'hDA;
            14'd8676: data_out = 8'hDE;
            14'd8677: data_out = 8'hFB;
            14'd8678: data_out = 8'hFD;
            14'd8679: data_out = 8'hFD;
            14'd8680: data_out = 8'hFD;
            14'd8681: data_out = 8'hFD;
            14'd8682: data_out = 8'hFD;
            14'd8683: data_out = 8'hFD;
            14'd8684: data_out = 8'hFD;
            14'd8685: data_out = 8'hFD;
            14'd8686: data_out = 8'hFC;
            14'd8687: data_out = 8'h7C;
            14'd8705: data_out = 8'h43;
            14'd8706: data_out = 8'h48;
            14'd8707: data_out = 8'hC8;
            14'd8708: data_out = 8'hFD;
            14'd8709: data_out = 8'hFD;
            14'd8710: data_out = 8'hFD;
            14'd8711: data_out = 8'hFD;
            14'd8712: data_out = 8'hFD;
            14'd8713: data_out = 8'hFD;
            14'd8714: data_out = 8'hFD;
            14'd8715: data_out = 8'hAF;
            14'd8735: data_out = 8'h78;
            14'd8736: data_out = 8'hFD;
            14'd8737: data_out = 8'hF9;
            14'd8738: data_out = 8'h98;
            14'd8739: data_out = 8'h33;
            14'd8740: data_out = 8'hA4;
            14'd8741: data_out = 8'hFD;
            14'd8742: data_out = 8'hFD;
            14'd8743: data_out = 8'hAF;
            14'd8763: data_out = 8'h32;
            14'd8764: data_out = 8'hFD;
            14'd8765: data_out = 8'hFD;
            14'd8766: data_out = 8'hFD;
            14'd8767: data_out = 8'hBC;
            14'd8768: data_out = 8'hFC;
            14'd8769: data_out = 8'hFD;
            14'd8770: data_out = 8'hFD;
            14'd8771: data_out = 8'h94;
            14'd8792: data_out = 8'hA7;
            14'd8793: data_out = 8'hFD;
            14'd8794: data_out = 8'hFD;
            14'd8795: data_out = 8'hFD;
            14'd8796: data_out = 8'hFD;
            14'd8797: data_out = 8'hFA;
            14'd8798: data_out = 8'hAF;
            14'd8799: data_out = 8'h0B;
            14'd8820: data_out = 8'h17;
            14'd8821: data_out = 8'hB4;
            14'd8822: data_out = 8'hE7;
            14'd8823: data_out = 8'hFD;
            14'd8824: data_out = 8'hDD;
            14'd8825: data_out = 8'h80;
            14'd8850: data_out = 8'h5D;
            14'd8851: data_out = 8'h95;
            14'd8852: data_out = 8'h16;
            14'd9425: data_out = 8'h24;
            14'd9426: data_out = 8'h38;
            14'd9427: data_out = 8'h89;
            14'd9428: data_out = 8'hC9;
            14'd9429: data_out = 8'hC7;
            14'd9430: data_out = 8'h5F;
            14'd9431: data_out = 8'h25;
            14'd9451: data_out = 8'h2D;
            14'd9452: data_out = 8'h98;
            14'd9453: data_out = 8'hEA;
            14'd9454: data_out = 8'hFE;
            14'd9455: data_out = 8'hFE;
            14'd9456: data_out = 8'hFE;
            14'd9457: data_out = 8'hFE;
            14'd9458: data_out = 8'hFE;
            14'd9459: data_out = 8'hFA;
            14'd9460: data_out = 8'hD3;
            14'd9461: data_out = 8'h97;
            14'd9477: data_out = 8'h2E;
            14'd9478: data_out = 8'h99;
            14'd9479: data_out = 8'hF0;
            14'd9480: data_out = 8'hFE;
            14'd9481: data_out = 8'hFE;
            14'd9482: data_out = 8'hE3;
            14'd9483: data_out = 8'hA6;
            14'd9484: data_out = 8'h85;
            14'd9485: data_out = 8'hFB;
            14'd9486: data_out = 8'hC8;
            14'd9487: data_out = 8'hFE;
            14'd9488: data_out = 8'hE5;
            14'd9489: data_out = 8'hE1;
            14'd9490: data_out = 8'h68;
            14'd9504: data_out = 8'h99;
            14'd9505: data_out = 8'hEA;
            14'd9506: data_out = 8'hFE;
            14'd9507: data_out = 8'hFE;
            14'd9508: data_out = 8'hBB;
            14'd9509: data_out = 8'h8E;
            14'd9513: data_out = 8'hBF;
            14'd9514: data_out = 8'h28;
            14'd9515: data_out = 8'hC6;
            14'd9516: data_out = 8'hF6;
            14'd9517: data_out = 8'hDF;
            14'd9518: data_out = 8'hFD;
            14'd9519: data_out = 8'h15;
            14'd9531: data_out = 8'h7E;
            14'd9532: data_out = 8'hFD;
            14'd9533: data_out = 8'hFE;
            14'd9534: data_out = 8'hE9;
            14'd9535: data_out = 8'h80;
            14'd9536: data_out = 8'h0B;
            14'd9541: data_out = 8'hD2;
            14'd9542: data_out = 8'h2B;
            14'd9543: data_out = 8'h46;
            14'd9544: data_out = 8'hFE;
            14'd9545: data_out = 8'hFE;
            14'd9546: data_out = 8'hFE;
            14'd9547: data_out = 8'h15;
            14'd9558: data_out = 8'h48;
            14'd9559: data_out = 8'hF3;
            14'd9560: data_out = 8'hFE;
            14'd9561: data_out = 8'hE4;
            14'd9562: data_out = 8'h36;
            14'd9568: data_out = 8'h20;
            14'd9569: data_out = 8'h74;
            14'd9570: data_out = 8'hE1;
            14'd9571: data_out = 8'hF2;
            14'd9572: data_out = 8'hFE;
            14'd9573: data_out = 8'hFF;
            14'd9574: data_out = 8'hA2;
            14'd9586: data_out = 8'h4B;
            14'd9587: data_out = 8'hF0;
            14'd9588: data_out = 8'hFE;
            14'd9589: data_out = 8'hDF;
            14'd9590: data_out = 8'h6D;
            14'd9591: data_out = 8'h8A;
            14'd9592: data_out = 8'hB2;
            14'd9593: data_out = 8'hB2;
            14'd9594: data_out = 8'hA9;
            14'd9595: data_out = 8'hD2;
            14'd9596: data_out = 8'hFB;
            14'd9597: data_out = 8'hE7;
            14'd9598: data_out = 8'hFE;
            14'd9599: data_out = 8'hFE;
            14'd9600: data_out = 8'hFE;
            14'd9601: data_out = 8'hE8;
            14'd9602: data_out = 8'h26;
            14'd9615: data_out = 8'hAF;
            14'd9616: data_out = 8'hF4;
            14'd9617: data_out = 8'hFD;
            14'd9618: data_out = 8'hFF;
            14'd9619: data_out = 8'hFE;
            14'd9620: data_out = 8'hFE;
            14'd9621: data_out = 8'hFB;
            14'd9622: data_out = 8'hFE;
            14'd9623: data_out = 8'hFE;
            14'd9624: data_out = 8'hFE;
            14'd9625: data_out = 8'hFE;
            14'd9626: data_out = 8'hFE;
            14'd9627: data_out = 8'hFC;
            14'd9628: data_out = 8'hAB;
            14'd9629: data_out = 8'h19;
            14'd9644: data_out = 8'h10;
            14'd9645: data_out = 8'h88;
            14'd9646: data_out = 8'hC3;
            14'd9647: data_out = 8'hB0;
            14'd9648: data_out = 8'h92;
            14'd9649: data_out = 8'h99;
            14'd9650: data_out = 8'hC8;
            14'd9651: data_out = 8'hFE;
            14'd9652: data_out = 8'hFE;
            14'd9653: data_out = 8'hFE;
            14'd9654: data_out = 8'hFE;
            14'd9655: data_out = 8'h96;
            14'd9656: data_out = 8'h10;
            14'd9678: data_out = 8'hA2;
            14'd9679: data_out = 8'hFE;
            14'd9680: data_out = 8'hFE;
            14'd9681: data_out = 8'hF1;
            14'd9682: data_out = 8'h63;
            14'd9705: data_out = 8'h76;
            14'd9706: data_out = 8'hFA;
            14'd9707: data_out = 8'hFE;
            14'd9708: data_out = 8'hFE;
            14'd9709: data_out = 8'h5A;
            14'd9732: data_out = 8'h64;
            14'd9733: data_out = 8'hF2;
            14'd9734: data_out = 8'hFE;
            14'd9735: data_out = 8'hFE;
            14'd9736: data_out = 8'hD3;
            14'd9759: data_out = 8'h36;
            14'd9760: data_out = 8'hF1;
            14'd9761: data_out = 8'hFE;
            14'd9762: data_out = 8'hFE;
            14'd9763: data_out = 8'hF2;
            14'd9764: data_out = 8'h3B;
            14'd9787: data_out = 8'h83;
            14'd9788: data_out = 8'hFE;
            14'd9789: data_out = 8'hFE;
            14'd9790: data_out = 8'hF4;
            14'd9791: data_out = 8'h40;
            14'd9814: data_out = 8'h0D;
            14'd9815: data_out = 8'hF9;
            14'd9816: data_out = 8'hFE;
            14'd9817: data_out = 8'hFE;
            14'd9818: data_out = 8'h98;
            14'd9841: data_out = 8'h0C;
            14'd9842: data_out = 8'hE4;
            14'd9843: data_out = 8'hFE;
            14'd9844: data_out = 8'hFE;
            14'd9845: data_out = 8'hD0;
            14'd9869: data_out = 8'h4E;
            14'd9870: data_out = 8'hFF;
            14'd9871: data_out = 8'hFE;
            14'd9872: data_out = 8'hFE;
            14'd9873: data_out = 8'h42;
            14'd9897: data_out = 8'hD1;
            14'd9898: data_out = 8'hFE;
            14'd9899: data_out = 8'hFE;
            14'd9900: data_out = 8'h89;
            14'd9925: data_out = 8'hE3;
            14'd9926: data_out = 8'hFF;
            14'd9927: data_out = 8'hE9;
            14'd9928: data_out = 8'h19;
            14'd9953: data_out = 8'h71;
            14'd9954: data_out = 8'hFF;
            14'd9955: data_out = 8'h6C;
            14'd10363: data_out = 8'h3D;
            14'd10365: data_out = 8'h2A;
            14'd10366: data_out = 8'h76;
            14'd10367: data_out = 8'hC1;
            14'd10368: data_out = 8'h76;
            14'd10369: data_out = 8'h76;
            14'd10370: data_out = 8'h3D;
            14'd10389: data_out = 8'h0E;
            14'd10390: data_out = 8'hB3;
            14'd10391: data_out = 8'hF5;
            14'd10392: data_out = 8'hEC;
            14'd10393: data_out = 8'hF2;
            14'd10394: data_out = 8'hFE;
            14'd10395: data_out = 8'hFE;
            14'd10396: data_out = 8'hFE;
            14'd10397: data_out = 8'hFE;
            14'd10398: data_out = 8'hF5;
            14'd10399: data_out = 8'hEB;
            14'd10400: data_out = 8'h54;
            14'd10417: data_out = 8'h97;
            14'd10418: data_out = 8'hFE;
            14'd10419: data_out = 8'hFE;
            14'd10420: data_out = 8'hFE;
            14'd10421: data_out = 8'hD5;
            14'd10422: data_out = 8'hC0;
            14'd10423: data_out = 8'hB2;
            14'd10424: data_out = 8'hB2;
            14'd10425: data_out = 8'hB4;
            14'd10426: data_out = 8'hFE;
            14'd10427: data_out = 8'hFE;
            14'd10428: data_out = 8'hF1;
            14'd10429: data_out = 8'h2E;
            14'd10444: data_out = 8'h2B;
            14'd10445: data_out = 8'hEB;
            14'd10446: data_out = 8'hFE;
            14'd10447: data_out = 8'hE2;
            14'd10448: data_out = 8'h40;
            14'd10449: data_out = 8'h1C;
            14'd10450: data_out = 8'h0C;
            14'd10454: data_out = 8'h80;
            14'd10455: data_out = 8'hFC;
            14'd10456: data_out = 8'hFF;
            14'd10457: data_out = 8'hAD;
            14'd10458: data_out = 8'h11;
            14'd10472: data_out = 8'h38;
            14'd10473: data_out = 8'hFE;
            14'd10474: data_out = 8'hFD;
            14'd10475: data_out = 8'h6B;
            14'd10483: data_out = 8'h86;
            14'd10484: data_out = 8'hFA;
            14'd10485: data_out = 8'hFE;
            14'd10486: data_out = 8'h4B;
            14'd10500: data_out = 8'h3F;
            14'd10501: data_out = 8'hFE;
            14'd10502: data_out = 8'h9E;
            14'd10512: data_out = 8'hDD;
            14'd10513: data_out = 8'hFE;
            14'd10514: data_out = 8'h9D;
            14'd10528: data_out = 8'hC2;
            14'd10529: data_out = 8'hFE;
            14'd10530: data_out = 8'h67;
            14'd10540: data_out = 8'h96;
            14'd10541: data_out = 8'hFE;
            14'd10542: data_out = 8'hD5;
            14'd10555: data_out = 8'h22;
            14'd10556: data_out = 8'hDC;
            14'd10557: data_out = 8'hEF;
            14'd10558: data_out = 8'h3A;
            14'd10568: data_out = 8'h54;
            14'd10569: data_out = 8'hFE;
            14'd10570: data_out = 8'hD5;
            14'd10583: data_out = 8'h7E;
            14'd10584: data_out = 8'hFE;
            14'd10585: data_out = 8'hAB;
            14'd10596: data_out = 8'h54;
            14'd10597: data_out = 8'hFE;
            14'd10598: data_out = 8'hD5;
            14'd10611: data_out = 8'hD6;
            14'd10612: data_out = 8'hEF;
            14'd10613: data_out = 8'h3C;
            14'd10624: data_out = 8'h54;
            14'd10625: data_out = 8'hFE;
            14'd10626: data_out = 8'hD5;
            14'd10639: data_out = 8'hD6;
            14'd10640: data_out = 8'hC7;
            14'd10652: data_out = 8'h54;
            14'd10653: data_out = 8'hFE;
            14'd10654: data_out = 8'hD5;
            14'd10666: data_out = 8'h0B;
            14'd10667: data_out = 8'hDB;
            14'd10668: data_out = 8'hC7;
            14'd10680: data_out = 8'h54;
            14'd10681: data_out = 8'hFE;
            14'd10682: data_out = 8'hD5;
            14'd10694: data_out = 8'h62;
            14'd10695: data_out = 8'hFE;
            14'd10696: data_out = 8'hC7;
            14'd10708: data_out = 8'hA2;
            14'd10709: data_out = 8'hFE;
            14'd10710: data_out = 8'hD1;
            14'd10722: data_out = 8'h62;
            14'd10723: data_out = 8'hFE;
            14'd10724: data_out = 8'hC7;
            14'd10735: data_out = 8'h33;
            14'd10736: data_out = 8'hEE;
            14'd10737: data_out = 8'hFE;
            14'd10738: data_out = 8'h4B;
            14'd10750: data_out = 8'h62;
            14'd10751: data_out = 8'hFE;
            14'd10752: data_out = 8'hC7;
            14'd10762: data_out = 8'h33;
            14'd10763: data_out = 8'hA5;
            14'd10764: data_out = 8'hFE;
            14'd10765: data_out = 8'hC3;
            14'd10778: data_out = 8'h42;
            14'd10779: data_out = 8'hF1;
            14'd10780: data_out = 8'hC7;
            14'd10790: data_out = 8'hA7;
            14'd10791: data_out = 8'hFE;
            14'd10792: data_out = 8'hE3;
            14'd10793: data_out = 8'h37;
            14'd10807: data_out = 8'hD6;
            14'd10808: data_out = 8'hD5;
            14'd10809: data_out = 8'h14;
            14'd10815: data_out = 8'h2E;
            14'd10816: data_out = 8'h98;
            14'd10817: data_out = 8'hCA;
            14'd10818: data_out = 8'hFE;
            14'd10819: data_out = 8'hFE;
            14'd10820: data_out = 8'h3F;
            14'd10835: data_out = 8'hD6;
            14'd10836: data_out = 8'hFE;
            14'd10837: data_out = 8'hCC;
            14'd10838: data_out = 8'hB4;
            14'd10839: data_out = 8'hB4;
            14'd10840: data_out = 8'hB4;
            14'd10841: data_out = 8'hB4;
            14'd10842: data_out = 8'hB4;
            14'd10843: data_out = 8'hEB;
            14'd10844: data_out = 8'hFE;
            14'd10845: data_out = 8'hFE;
            14'd10846: data_out = 8'hEA;
            14'd10847: data_out = 8'h9C;
            14'd10863: data_out = 8'h51;
            14'd10864: data_out = 8'hCD;
            14'd10865: data_out = 8'hFE;
            14'd10866: data_out = 8'hFE;
            14'd10867: data_out = 8'hFE;
            14'd10868: data_out = 8'hFE;
            14'd10869: data_out = 8'hFE;
            14'd10870: data_out = 8'hFE;
            14'd10871: data_out = 8'hFE;
            14'd10872: data_out = 8'hFC;
            14'd10873: data_out = 8'hEA;
            14'd10874: data_out = 8'h78;
            14'd10892: data_out = 8'h1A;
            14'd10893: data_out = 8'hD2;
            14'd10894: data_out = 8'hFE;
            14'd10895: data_out = 8'hFE;
            14'd10896: data_out = 8'hFE;
            14'd10897: data_out = 8'hFE;
            14'd10898: data_out = 8'hFE;
            14'd10899: data_out = 8'h99;
            14'd10900: data_out = 8'h68;
            14'd11359: data_out = 8'hCC;
            14'd11360: data_out = 8'hFD;
            14'd11361: data_out = 8'hB0;
            14'd11386: data_out = 8'h96;
            14'd11387: data_out = 8'hFC;
            14'd11388: data_out = 8'hFC;
            14'd11389: data_out = 8'h7D;
            14'd11413: data_out = 8'h75;
            14'd11414: data_out = 8'hFC;
            14'd11415: data_out = 8'hBA;
            14'd11416: data_out = 8'h38;
            14'd11441: data_out = 8'h8D;
            14'd11442: data_out = 8'hFC;
            14'd11443: data_out = 8'h76;
            14'd11469: data_out = 8'h9A;
            14'd11470: data_out = 8'hF7;
            14'd11471: data_out = 8'h32;
            14'd11496: data_out = 8'h1A;
            14'd11497: data_out = 8'hFD;
            14'd11498: data_out = 8'hC4;
            14'd11524: data_out = 8'h96;
            14'd11525: data_out = 8'hFD;
            14'd11526: data_out = 8'hC4;
            14'd11534: data_out = 8'h39;
            14'd11535: data_out = 8'h55;
            14'd11536: data_out = 8'h55;
            14'd11537: data_out = 8'h26;
            14'd11552: data_out = 8'hE1;
            14'd11553: data_out = 8'hFD;
            14'd11554: data_out = 8'h60;
            14'd11560: data_out = 8'h97;
            14'd11561: data_out = 8'hE2;
            14'd11562: data_out = 8'hF3;
            14'd11563: data_out = 8'hFC;
            14'd11564: data_out = 8'hFC;
            14'd11565: data_out = 8'hEE;
            14'd11566: data_out = 8'h7D;
            14'd11580: data_out = 8'hE5;
            14'd11581: data_out = 8'hE2;
            14'd11586: data_out = 8'h36;
            14'd11587: data_out = 8'hE5;
            14'd11588: data_out = 8'hFD;
            14'd11589: data_out = 8'hFF;
            14'd11590: data_out = 8'hEA;
            14'd11591: data_out = 8'hAF;
            14'd11592: data_out = 8'hE1;
            14'd11593: data_out = 8'hFF;
            14'd11594: data_out = 8'hE4;
            14'd11595: data_out = 8'h1F;
            14'd11607: data_out = 8'h6E;
            14'd11608: data_out = 8'hFC;
            14'd11609: data_out = 8'h96;
            14'd11612: data_out = 8'h1A;
            14'd11613: data_out = 8'h80;
            14'd11614: data_out = 8'hFC;
            14'd11615: data_out = 8'hFC;
            14'd11616: data_out = 8'hE3;
            14'd11617: data_out = 8'h86;
            14'd11618: data_out = 8'h1C;
            14'd11621: data_out = 8'hB2;
            14'd11622: data_out = 8'hFC;
            14'd11623: data_out = 8'h38;
            14'd11635: data_out = 8'h9F;
            14'd11636: data_out = 8'hFC;
            14'd11637: data_out = 8'h71;
            14'd11640: data_out = 8'h96;
            14'd11641: data_out = 8'hFD;
            14'd11642: data_out = 8'hFC;
            14'd11643: data_out = 8'hBA;
            14'd11644: data_out = 8'h2B;
            14'd11649: data_out = 8'h8D;
            14'd11650: data_out = 8'hFC;
            14'd11651: data_out = 8'h38;
            14'd11663: data_out = 8'hB9;
            14'd11664: data_out = 8'hFC;
            14'd11665: data_out = 8'h71;
            14'd11667: data_out = 8'h26;
            14'd11668: data_out = 8'hED;
            14'd11669: data_out = 8'hFD;
            14'd11670: data_out = 8'h97;
            14'd11677: data_out = 8'h8D;
            14'd11678: data_out = 8'hCA;
            14'd11691: data_out = 8'hC6;
            14'd11692: data_out = 8'hFD;
            14'd11693: data_out = 8'h72;
            14'd11695: data_out = 8'h93;
            14'd11696: data_out = 8'hFD;
            14'd11697: data_out = 8'hA3;
            14'd11705: data_out = 8'h9A;
            14'd11706: data_out = 8'hC5;
            14'd11719: data_out = 8'hC5;
            14'd11720: data_out = 8'hFC;
            14'd11721: data_out = 8'h71;
            14'd11723: data_out = 8'hAC;
            14'd11724: data_out = 8'hFC;
            14'd11725: data_out = 8'hBC;
            14'd11732: data_out = 8'h1A;
            14'd11733: data_out = 8'hFD;
            14'd11734: data_out = 8'hAB;
            14'd11747: data_out = 8'hC5;
            14'd11748: data_out = 8'hFC;
            14'd11749: data_out = 8'h71;
            14'd11751: data_out = 8'h13;
            14'd11752: data_out = 8'hE7;
            14'd11753: data_out = 8'hF7;
            14'd11754: data_out = 8'h7A;
            14'd11755: data_out = 8'h13;
            14'd11760: data_out = 8'hC8;
            14'd11761: data_out = 8'hF4;
            14'd11762: data_out = 8'h38;
            14'd11774: data_out = 8'h1A;
            14'd11775: data_out = 8'hDE;
            14'd11776: data_out = 8'hFC;
            14'd11777: data_out = 8'h71;
            14'd11780: data_out = 8'h19;
            14'd11781: data_out = 8'hCB;
            14'd11782: data_out = 8'hFC;
            14'd11783: data_out = 8'hC1;
            14'd11784: data_out = 8'h0D;
            14'd11786: data_out = 8'h4C;
            14'd11787: data_out = 8'hC8;
            14'd11788: data_out = 8'hF9;
            14'd11789: data_out = 8'h7D;
            14'd11803: data_out = 8'hB9;
            14'd11804: data_out = 8'hFD;
            14'd11805: data_out = 8'hB3;
            14'd11810: data_out = 8'h4C;
            14'd11811: data_out = 8'h23;
            14'd11812: data_out = 8'h1D;
            14'd11813: data_out = 8'h9A;
            14'd11814: data_out = 8'hFD;
            14'd11815: data_out = 8'hF4;
            14'd11816: data_out = 8'h7D;
            14'd11831: data_out = 8'h1C;
            14'd11832: data_out = 8'hD1;
            14'd11833: data_out = 8'hFD;
            14'd11834: data_out = 8'hC4;
            14'd11835: data_out = 8'h52;
            14'd11836: data_out = 8'h39;
            14'd11837: data_out = 8'h39;
            14'd11838: data_out = 8'h83;
            14'd11839: data_out = 8'hC5;
            14'd11840: data_out = 8'hFC;
            14'd11841: data_out = 8'hFD;
            14'd11842: data_out = 8'hD6;
            14'd11843: data_out = 8'h51;
            14'd11860: data_out = 8'h19;
            14'd11861: data_out = 8'hD8;
            14'd11862: data_out = 8'hFC;
            14'd11863: data_out = 8'hFC;
            14'd11864: data_out = 8'hFC;
            14'd11865: data_out = 8'hFD;
            14'd11866: data_out = 8'hFC;
            14'd11867: data_out = 8'hFC;
            14'd11868: data_out = 8'hFC;
            14'd11869: data_out = 8'h9C;
            14'd11870: data_out = 8'h13;
            14'd11889: data_out = 8'h10;
            14'd11890: data_out = 8'h67;
            14'd11891: data_out = 8'h8B;
            14'd11892: data_out = 8'hF0;
            14'd11893: data_out = 8'h8C;
            14'd11894: data_out = 8'h8B;
            14'd11895: data_out = 8'h8B;
            14'd11896: data_out = 8'h28;
            14'd12496: data_out = 8'h31;
            14'd12497: data_out = 8'hB4;
            14'd12498: data_out = 8'hFD;
            14'd12499: data_out = 8'hFF;
            14'd12500: data_out = 8'hFD;
            14'd12501: data_out = 8'hA9;
            14'd12502: data_out = 8'h24;
            14'd12503: data_out = 8'h0B;
            14'd12504: data_out = 8'h4C;
            14'd12523: data_out = 8'h44;
            14'd12524: data_out = 8'hE4;
            14'd12525: data_out = 8'hFC;
            14'd12526: data_out = 8'hFC;
            14'd12527: data_out = 8'hFD;
            14'd12528: data_out = 8'hFC;
            14'd12529: data_out = 8'hFC;
            14'd12530: data_out = 8'hA0;
            14'd12531: data_out = 8'hBD;
            14'd12532: data_out = 8'hFD;
            14'd12533: data_out = 8'h5C;
            14'd12550: data_out = 8'h37;
            14'd12551: data_out = 8'hFC;
            14'd12552: data_out = 8'hFC;
            14'd12553: data_out = 8'hE3;
            14'd12554: data_out = 8'h4F;
            14'd12555: data_out = 8'h45;
            14'd12556: data_out = 8'h45;
            14'd12557: data_out = 8'h64;
            14'd12558: data_out = 8'h5A;
            14'd12559: data_out = 8'hEC;
            14'd12560: data_out = 8'hF7;
            14'd12561: data_out = 8'h43;
            14'd12577: data_out = 8'h2B;
            14'd12578: data_out = 8'hE9;
            14'd12579: data_out = 8'hFC;
            14'd12580: data_out = 8'hB9;
            14'd12581: data_out = 8'h32;
            14'd12585: data_out = 8'h1A;
            14'd12586: data_out = 8'hCB;
            14'd12587: data_out = 8'hFC;
            14'd12588: data_out = 8'h87;
            14'd12605: data_out = 8'hA8;
            14'd12606: data_out = 8'hFD;
            14'd12607: data_out = 8'hB2;
            14'd12608: data_out = 8'h25;
            14'd12613: data_out = 8'h46;
            14'd12614: data_out = 8'hFC;
            14'd12615: data_out = 8'hFC;
            14'd12616: data_out = 8'h3F;
            14'd12632: data_out = 8'h9B;
            14'd12633: data_out = 8'hFD;
            14'd12634: data_out = 8'hF2;
            14'd12635: data_out = 8'h2A;
            14'd12641: data_out = 8'hBF;
            14'd12642: data_out = 8'hFD;
            14'd12643: data_out = 8'hBE;
            14'd12660: data_out = 8'hCF;
            14'd12661: data_out = 8'hFC;
            14'd12662: data_out = 8'hE6;
            14'd12668: data_out = 8'h88;
            14'd12669: data_out = 8'hFC;
            14'd12670: data_out = 8'hFC;
            14'd12671: data_out = 8'h40;
            14'd12688: data_out = 8'hCF;
            14'd12689: data_out = 8'hFC;
            14'd12690: data_out = 8'hE6;
            14'd12694: data_out = 8'h20;
            14'd12695: data_out = 8'h8A;
            14'd12696: data_out = 8'hFC;
            14'd12697: data_out = 8'hFC;
            14'd12698: data_out = 8'hE3;
            14'd12699: data_out = 8'h10;
            14'd12716: data_out = 8'hA5;
            14'd12717: data_out = 8'hFC;
            14'd12718: data_out = 8'hF9;
            14'd12719: data_out = 8'hCF;
            14'd12720: data_out = 8'hCF;
            14'd12721: data_out = 8'hCF;
            14'd12722: data_out = 8'hE4;
            14'd12723: data_out = 8'hFD;
            14'd12724: data_out = 8'hFC;
            14'd12725: data_out = 8'hFC;
            14'd12726: data_out = 8'hA0;
            14'd12745: data_out = 8'hB3;
            14'd12746: data_out = 8'hFD;
            14'd12747: data_out = 8'hFC;
            14'd12748: data_out = 8'hFC;
            14'd12749: data_out = 8'hFC;
            14'd12750: data_out = 8'hFC;
            14'd12751: data_out = 8'h4B;
            14'd12752: data_out = 8'hA9;
            14'd12753: data_out = 8'hFC;
            14'd12754: data_out = 8'h38;
            14'd12774: data_out = 8'h40;
            14'd12775: data_out = 8'h74;
            14'd12776: data_out = 8'h74;
            14'd12777: data_out = 8'h4A;
            14'd12779: data_out = 8'h95;
            14'd12780: data_out = 8'hFD;
            14'd12781: data_out = 8'hD7;
            14'd12782: data_out = 8'h15;
            14'd12807: data_out = 8'hFD;
            14'd12808: data_out = 8'hFC;
            14'd12809: data_out = 8'hA2;
            14'd12834: data_out = 8'h20;
            14'd12835: data_out = 8'hFD;
            14'd12836: data_out = 8'hF0;
            14'd12837: data_out = 8'h32;
            14'd12862: data_out = 8'h9D;
            14'd12863: data_out = 8'hFD;
            14'd12864: data_out = 8'hA4;
            14'd12889: data_out = 8'h2B;
            14'd12890: data_out = 8'hF0;
            14'd12891: data_out = 8'hFD;
            14'd12892: data_out = 8'h5C;
            14'd12917: data_out = 8'h5D;
            14'd12918: data_out = 8'hFD;
            14'd12919: data_out = 8'hFC;
            14'd12920: data_out = 8'h54;
            14'd12945: data_out = 8'h72;
            14'd12946: data_out = 8'hFC;
            14'd12947: data_out = 8'hD1;
            14'd12973: data_out = 8'hCF;
            14'd12974: data_out = 8'hFC;
            14'd12975: data_out = 8'h74;
            14'd13001: data_out = 8'hA5;
            14'd13002: data_out = 8'hFC;
            14'd13003: data_out = 8'h74;
            14'd13029: data_out = 8'h5D;
            14'd13030: data_out = 8'hC8;
            14'd13031: data_out = 8'h3F;
            14'd13464: data_out = 8'h11;
            14'd13465: data_out = 8'h42;
            14'd13466: data_out = 8'h8A;
            14'd13467: data_out = 8'hFF;
            14'd13468: data_out = 8'hFD;
            14'd13469: data_out = 8'hA9;
            14'd13470: data_out = 8'h8A;
            14'd13471: data_out = 8'h17;
            14'd13491: data_out = 8'h78;
            14'd13492: data_out = 8'hE4;
            14'd13493: data_out = 8'hFC;
            14'd13494: data_out = 8'hFC;
            14'd13495: data_out = 8'hFD;
            14'd13496: data_out = 8'hFC;
            14'd13497: data_out = 8'hFC;
            14'd13498: data_out = 8'hFC;
            14'd13499: data_out = 8'h9E;
            14'd13518: data_out = 8'h6C;
            14'd13519: data_out = 8'hFC;
            14'd13520: data_out = 8'hFC;
            14'd13521: data_out = 8'hFC;
            14'd13522: data_out = 8'hFC;
            14'd13523: data_out = 8'hBE;
            14'd13524: data_out = 8'hFC;
            14'd13525: data_out = 8'hFC;
            14'd13526: data_out = 8'hFC;
            14'd13527: data_out = 8'hFC;
            14'd13545: data_out = 8'h2B;
            14'd13546: data_out = 8'hE9;
            14'd13547: data_out = 8'hFC;
            14'd13548: data_out = 8'hFC;
            14'd13549: data_out = 8'hFC;
            14'd13550: data_out = 8'h74;
            14'd13552: data_out = 8'h87;
            14'd13553: data_out = 8'hFC;
            14'd13554: data_out = 8'hFC;
            14'd13555: data_out = 8'hFC;
            14'd13572: data_out = 8'h2B;
            14'd13573: data_out = 8'hB2;
            14'd13574: data_out = 8'hFD;
            14'd13575: data_out = 8'hFC;
            14'd13576: data_out = 8'hDD;
            14'd13577: data_out = 8'h2B;
            14'd13581: data_out = 8'h36;
            14'd13582: data_out = 8'hE8;
            14'd13583: data_out = 8'hFC;
            14'd13584: data_out = 8'hD2;
            14'd13600: data_out = 8'h5D;
            14'd13601: data_out = 8'hFD;
            14'd13602: data_out = 8'hFF;
            14'd13603: data_out = 8'hF9;
            14'd13604: data_out = 8'h73;
            14'd13610: data_out = 8'h88;
            14'd13611: data_out = 8'hFB;
            14'd13612: data_out = 8'hFF;
            14'd13613: data_out = 8'h9A;
            14'd13628: data_out = 8'hA6;
            14'd13629: data_out = 8'hFC;
            14'd13630: data_out = 8'hFD;
            14'd13631: data_out = 8'hB9;
            14'd13639: data_out = 8'hD1;
            14'd13640: data_out = 8'hFD;
            14'd13641: data_out = 8'hCE;
            14'd13655: data_out = 8'h13;
            14'd13656: data_out = 8'hDC;
            14'd13657: data_out = 8'hFC;
            14'd13658: data_out = 8'hFD;
            14'd13659: data_out = 8'h5C;
            14'd13667: data_out = 8'h74;
            14'd13668: data_out = 8'hFD;
            14'd13669: data_out = 8'hCE;
            14'd13683: data_out = 8'h46;
            14'd13684: data_out = 8'hFC;
            14'd13685: data_out = 8'hFC;
            14'd13686: data_out = 8'hC0;
            14'd13687: data_out = 8'h11;
            14'd13695: data_out = 8'h74;
            14'd13696: data_out = 8'hFD;
            14'd13697: data_out = 8'hDF;
            14'd13698: data_out = 8'h19;
            14'd13711: data_out = 8'h7A;
            14'd13712: data_out = 8'hFC;
            14'd13713: data_out = 8'hFC;
            14'd13714: data_out = 8'h3F;
            14'd13723: data_out = 8'h74;
            14'd13724: data_out = 8'hFD;
            14'd13725: data_out = 8'hFC;
            14'd13726: data_out = 8'h45;
            14'd13739: data_out = 8'h84;
            14'd13740: data_out = 8'hFD;
            14'd13741: data_out = 8'hFD;
            14'd13751: data_out = 8'h74;
            14'd13752: data_out = 8'hFF;
            14'd13753: data_out = 8'hFD;
            14'd13754: data_out = 8'h45;
            14'd13767: data_out = 8'hB8;
            14'd13768: data_out = 8'hFC;
            14'd13769: data_out = 8'hFC;
            14'd13779: data_out = 8'h74;
            14'd13780: data_out = 8'hFD;
            14'd13781: data_out = 8'hFC;
            14'd13782: data_out = 8'h45;
            14'd13795: data_out = 8'hB8;
            14'd13796: data_out = 8'hFC;
            14'd13797: data_out = 8'hFC;
            14'd13807: data_out = 8'h74;
            14'd13808: data_out = 8'hFD;
            14'd13809: data_out = 8'hF0;
            14'd13810: data_out = 8'h32;
            14'd13823: data_out = 8'hB8;
            14'd13824: data_out = 8'hFC;
            14'd13825: data_out = 8'hFC;
            14'd13835: data_out = 8'hD2;
            14'd13836: data_out = 8'hFD;
            14'd13837: data_out = 8'h70;
            14'd13851: data_out = 8'h30;
            14'd13852: data_out = 8'hE8;
            14'd13853: data_out = 8'hFC;
            14'd13854: data_out = 8'h9E;
            14'd13863: data_out = 8'hE6;
            14'd13864: data_out = 8'hE8;
            14'd13880: data_out = 8'h5D;
            14'd13881: data_out = 8'hFD;
            14'd13882: data_out = 8'hF4;
            14'd13883: data_out = 8'h32;
            14'd13890: data_out = 8'h9B;
            14'd13891: data_out = 8'hFD;
            14'd13892: data_out = 8'hA8;
            14'd13908: data_out = 8'h22;
            14'd13909: data_out = 8'hA4;
            14'd13910: data_out = 8'hFD;
            14'd13911: data_out = 8'h71;
            14'd13917: data_out = 8'h42;
            14'd13918: data_out = 8'hEC;
            14'd13919: data_out = 8'hE7;
            14'd13920: data_out = 8'h2A;
            14'd13937: data_out = 8'h20;
            14'd13938: data_out = 8'hDE;
            14'd13939: data_out = 8'hF0;
            14'd13940: data_out = 8'h86;
            14'd13943: data_out = 8'h26;
            14'd13944: data_out = 8'h5B;
            14'd13945: data_out = 8'hEA;
            14'd13946: data_out = 8'hFC;
            14'd13947: data_out = 8'h89;
            14'd13966: data_out = 8'h19;
            14'd13967: data_out = 8'hB1;
            14'd13968: data_out = 8'hF0;
            14'd13969: data_out = 8'hCF;
            14'd13970: data_out = 8'h67;
            14'd13971: data_out = 8'hE9;
            14'd13972: data_out = 8'hFC;
            14'd13973: data_out = 8'hFC;
            14'd13974: data_out = 8'hB0;
            14'd13975: data_out = 8'h23;
            14'd13995: data_out = 8'h0F;
            14'd13996: data_out = 8'h36;
            14'd13997: data_out = 8'hB3;
            14'd13998: data_out = 8'hFC;
            14'd13999: data_out = 8'h89;
            14'd14000: data_out = 8'h89;
            14'd14001: data_out = 8'h36;
            14'd14461: data_out = 8'h80;
            14'd14462: data_out = 8'hFF;
            14'd14463: data_out = 8'hBF;
            14'd14489: data_out = 8'hBF;
            14'd14490: data_out = 8'hFF;
            14'd14491: data_out = 8'hFF;
            14'd14492: data_out = 8'h40;
            14'd14517: data_out = 8'hFF;
            14'd14518: data_out = 8'hFF;
            14'd14519: data_out = 8'hFF;
            14'd14520: data_out = 8'h80;
            14'd14545: data_out = 8'hFF;
            14'd14546: data_out = 8'hFF;
            14'd14547: data_out = 8'hFF;
            14'd14573: data_out = 8'hFF;
            14'd14574: data_out = 8'hFF;
            14'd14575: data_out = 8'hFF;
            14'd14601: data_out = 8'h80;
            14'd14602: data_out = 8'hFF;
            14'd14603: data_out = 8'hFF;
            14'd14604: data_out = 8'h80;
            14'd14629: data_out = 8'hFF;
            14'd14630: data_out = 8'hFF;
            14'd14631: data_out = 8'hFF;
            14'd14632: data_out = 8'h80;
            14'd14657: data_out = 8'hFF;
            14'd14658: data_out = 8'hFF;
            14'd14659: data_out = 8'hFF;
            14'd14660: data_out = 8'h80;
            14'd14685: data_out = 8'hFF;
            14'd14686: data_out = 8'hFF;
            14'd14687: data_out = 8'hFF;
            14'd14688: data_out = 8'h80;
            14'd14713: data_out = 8'hFF;
            14'd14714: data_out = 8'hFF;
            14'd14715: data_out = 8'hFF;
            14'd14716: data_out = 8'h80;
            14'd14741: data_out = 8'hFF;
            14'd14742: data_out = 8'hFF;
            14'd14743: data_out = 8'hFF;
            14'd14769: data_out = 8'hFF;
            14'd14770: data_out = 8'hFF;
            14'd14771: data_out = 8'hFF;
            14'd14797: data_out = 8'hFF;
            14'd14798: data_out = 8'hFF;
            14'd14799: data_out = 8'hFF;
            14'd14825: data_out = 8'hFF;
            14'd14826: data_out = 8'hFF;
            14'd14827: data_out = 8'hFF;
            14'd14853: data_out = 8'hBF;
            14'd14854: data_out = 8'hFF;
            14'd14855: data_out = 8'hFF;
            14'd14856: data_out = 8'h80;
            14'd14881: data_out = 8'hBF;
            14'd14882: data_out = 8'hFF;
            14'd14883: data_out = 8'hFF;
            14'd14884: data_out = 8'h80;
            14'd14908: data_out = 8'h40;
            14'd14909: data_out = 8'hFF;
            14'd14910: data_out = 8'hFF;
            14'd14911: data_out = 8'hFF;
            14'd14912: data_out = 8'h80;
            14'd14936: data_out = 8'hBF;
            14'd14937: data_out = 8'hFF;
            14'd14938: data_out = 8'hFF;
            14'd14939: data_out = 8'hFF;
            14'd14940: data_out = 8'h80;
            14'd14963: data_out = 8'h40;
            14'd14964: data_out = 8'hFF;
            14'd14965: data_out = 8'hFF;
            14'd14966: data_out = 8'hFF;
            14'd14967: data_out = 8'h40;
            14'd14991: data_out = 8'h40;
            14'd14992: data_out = 8'hFF;
            14'd14993: data_out = 8'h80;
            14'd15484: data_out = 8'h33;
            14'd15485: data_out = 8'h84;
            14'd15486: data_out = 8'hD6;
            14'd15487: data_out = 8'hFD;
            14'd15488: data_out = 8'hFE;
            14'd15489: data_out = 8'hFD;
            14'd15490: data_out = 8'hCB;
            14'd15491: data_out = 8'hA2;
            14'd15492: data_out = 8'h29;
            14'd15508: data_out = 8'h66;
            14'd15509: data_out = 8'h8E;
            14'd15510: data_out = 8'hCB;
            14'd15511: data_out = 8'hCB;
            14'd15512: data_out = 8'hFD;
            14'd15513: data_out = 8'hFC;
            14'd15514: data_out = 8'hFD;
            14'd15515: data_out = 8'hFC;
            14'd15516: data_out = 8'h97;
            14'd15517: data_out = 8'h46;
            14'd15536: data_out = 8'hFE;
            14'd15537: data_out = 8'hFD;
            14'd15538: data_out = 8'hF4;
            14'd15539: data_out = 8'hCB;
            14'd15540: data_out = 8'h8E;
            14'd15541: data_out = 8'h66;
            14'd15542: data_out = 8'h52;
            14'd15564: data_out = 8'hAC;
            14'd15565: data_out = 8'hFC;
            14'd15566: data_out = 8'hCB;
            14'd15592: data_out = 8'h15;
            14'd15593: data_out = 8'hDF;
            14'd15594: data_out = 8'hEA;
            14'd15595: data_out = 8'h1E;
            14'd15621: data_out = 8'h7A;
            14'd15622: data_out = 8'hFD;
            14'd15623: data_out = 8'h32;
            14'd15649: data_out = 8'h7B;
            14'd15650: data_out = 8'hFE;
            14'd15651: data_out = 8'h5B;
            14'd15652: data_out = 8'h33;
            14'd15653: data_out = 8'h33;
            14'd15654: data_out = 8'h33;
            14'd15676: data_out = 8'h15;
            14'd15677: data_out = 8'hDF;
            14'd15678: data_out = 8'hFD;
            14'd15679: data_out = 8'hFC;
            14'd15680: data_out = 8'hFD;
            14'd15681: data_out = 8'hFC;
            14'd15682: data_out = 8'hFD;
            14'd15683: data_out = 8'hAC;
            14'd15684: data_out = 8'h52;
            14'd15703: data_out = 8'h15;
            14'd15704: data_out = 8'hD6;
            14'd15705: data_out = 8'hFD;
            14'd15706: data_out = 8'hCB;
            14'd15707: data_out = 8'hA2;
            14'd15708: data_out = 8'h66;
            14'd15709: data_out = 8'h66;
            14'd15710: data_out = 8'hCB;
            14'd15711: data_out = 8'hDF;
            14'd15712: data_out = 8'hFE;
            14'd15713: data_out = 8'hFD;
            14'd15714: data_out = 8'h33;
            14'd15731: data_out = 8'h3D;
            14'd15732: data_out = 8'hFD;
            14'd15733: data_out = 8'hAB;
            14'd15739: data_out = 8'h14;
            14'd15740: data_out = 8'h70;
            14'd15741: data_out = 8'hC0;
            14'd15742: data_out = 8'hFD;
            14'd15743: data_out = 8'hD4;
            14'd15744: data_out = 8'h29;
            14'd15770: data_out = 8'h66;
            14'd15771: data_out = 8'hCB;
            14'd15772: data_out = 8'hEA;
            14'd15773: data_out = 8'h33;
            14'd15799: data_out = 8'h14;
            14'd15800: data_out = 8'hD5;
            14'd15801: data_out = 8'hE8;
            14'd15802: data_out = 8'h52;
            14'd15828: data_out = 8'h3E;
            14'd15829: data_out = 8'hCB;
            14'd15830: data_out = 8'hEA;
            14'd15831: data_out = 8'h70;
            14'd15857: data_out = 8'h14;
            14'd15858: data_out = 8'hD5;
            14'd15859: data_out = 8'hFC;
            14'd15886: data_out = 8'h99;
            14'd15887: data_out = 8'hFD;
            14'd15913: data_out = 8'h29;
            14'd15914: data_out = 8'hE9;
            14'd15915: data_out = 8'hD4;
            14'd15928: data_out = 8'h71;
            14'd15929: data_out = 8'h5C;
            14'd15940: data_out = 8'h1F;
            14'd15941: data_out = 8'hAD;
            14'd15942: data_out = 8'hF4;
            14'd15943: data_out = 8'h28;
            14'd15955: data_out = 8'h52;
            14'd15956: data_out = 8'hFD;
            14'd15957: data_out = 8'h97;
            14'd15964: data_out = 8'h15;
            14'd15965: data_out = 8'h66;
            14'd15966: data_out = 8'h66;
            14'd15967: data_out = 8'hB7;
            14'd15968: data_out = 8'hE9;
            14'd15969: data_out = 8'hD4;
            14'd15970: data_out = 8'h51;
            14'd15983: data_out = 8'h52;
            14'd15984: data_out = 8'hFF;
            14'd15985: data_out = 8'hFD;
            14'd15986: data_out = 8'hEA;
            14'd15987: data_out = 8'h98;
            14'd15988: data_out = 8'h99;
            14'd15989: data_out = 8'hC1;
            14'd15990: data_out = 8'hAD;
            14'd15991: data_out = 8'hFD;
            14'd15992: data_out = 8'hFE;
            14'd15993: data_out = 8'hFD;
            14'd15994: data_out = 8'hFE;
            14'd15995: data_out = 8'hD5;
            14'd15996: data_out = 8'h8E;
            14'd15997: data_out = 8'h14;
            14'd16012: data_out = 8'h47;
            14'd16013: data_out = 8'h97;
            14'd16014: data_out = 8'h97;
            14'd16015: data_out = 8'hE8;
            14'd16016: data_out = 8'hFD;
            14'd16017: data_out = 8'hD4;
            14'd16018: data_out = 8'hC0;
            14'd16019: data_out = 8'h97;
            14'd16020: data_out = 8'h83;
            14'd16021: data_out = 8'h32;
            14'd16022: data_out = 8'h32;
            default: data_out = 8'h00;
        endcase
    end
endmodule
