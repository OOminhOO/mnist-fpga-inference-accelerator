`timescale 1ns / 1ps

module tb_cnn_1k_verify;

    // ========================================================================
    // 1. �Ķ���� �� ��� ���� (�ڼ��� �ʿ��)
    // ========================================================================
    // �Ʊ� �����Ͻ� ���� ��η� �����ּ���!
    parameter IMG_FILE = "input_1k.txt";
    parameter LBL_FILE = "label_1k.txt";

    integer N_TEST = 1000; // �׽�Ʈ�� ����

    // ========================================================================
    // 2. ��ȣ ����
    // ========================================================================
    reg          clk;
    reg          rst_n;
    reg  [7:0]   data_in;
    reg          data_valid;
    wire [3:0]   decision;
    wire         out_valid;

    // ��뷮 �޸� ����
    // 1000�� * 784�ȼ� = 784,000 ����Ʈ
    reg [7:0]  mem_inputs [0:784000]; 
    reg [31:0] mem_labels [0:1000];   // ������

    // ī���� �� �ε���
    integer img_idx;   // �� ��° �̹�������
    integer px_idx;    // �ȼ� �ε��� (0~783)
    integer correct_cnt;
    integer error_cnt;
    integer file_ptr_idx; // ��ü �޸� �ε���

    // ========================================================================
    // 3. DUT �ν��Ͻ�
    // ========================================================================
    cnn_core_top u_dut (
        .clk        (clk),
        .rst_n      (rst_n),
        .data_in    (data_in),
        .data_valid (data_valid),
        .decision   (decision),
        .out_valid  (out_valid)
    );

    // ========================================================================
    // 4. Ŭ�� �� �ʱ�ȭ
    // ========================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 100MHz
    end

    // ========================================================================
    // 5. ���� ���� ������
    // ========================================================================
    initial begin
        // (1) ���� �ε�
        $display("\n[TB] Loading 1,000 Images & Labels...");
        $readmemh(IMG_FILE, mem_inputs);
        $readmemh(LBL_FILE, mem_labels);

        // (2) ���� �ʱ�ȭ
        rst_n = 0;
        data_valid = 0;
        data_in = 0;
        correct_cnt = 0;
        error_cnt = 0;
        
        #100;
        rst_n = 1;
        #100;

        $display("[TB] Start 1,000 Image Verification Loop...");
        $display("------------------------------------------------");

        // (3) ���� ����
        for (img_idx = 0; img_idx < N_TEST; img_idx = img_idx + 1) begin
            
            // --- �̹��� 1�� ���� (784Ŭ��) ---
            for (px_idx = 0; px_idx < 784; px_idx = px_idx + 1) begin
                @(posedge clk);
                data_valid <= 1;
                // �޸� �ּ� ���: (���� �̹��� ��ȣ * 784) + �ȼ� ��ȣ
                data_in    <= mem_inputs[img_idx * 784 + px_idx];
            end
            
            // ���� ��
            @(posedge clk);
            data_valid <= 0;
            data_in    <= 0;

            // --- ��� ��� ---
            // out_valid�� 1�� �� ������ ��ٸ�
            wait(out_valid);
            
            // --- ä�� ---
            // Ÿ�̹� ���߱� ���� Ŭ�� �������� ���ø�
            @(posedge clk); 
            if (decision === mem_labels[img_idx][3:0]) begin
                correct_cnt = correct_cnt + 1;
            end else begin
                error_cnt = error_cnt + 1;
                $display("[FAIL] Image #%0d: Expected=%d, Got=%d", 
                         img_idx, mem_labels[img_idx], decision);
            end

            // ���� ��Ȳ ��� (100������)
            if ((img_idx + 1) % 100 == 0) begin
                $display("   ... Processed %0d/%0d (Errors: %0d)", 
                         img_idx + 1, N_TEST, error_cnt);
            end

            // ���� �̹����� ���� �ణ�� ���� �� (Pipeline Flush ����)
            repeat(20) @(posedge clk);
        end

        // (4) ���� ��� ���
        $display("------------------------------------------------");
        $display("[FINAL RESULT]");
        $display("Total Images : %0d", N_TEST);
        $display("Correct      : %0d", correct_cnt);
        $display("Errors       : %0d", error_cnt);
        
        if (error_cnt == 0) begin
            $display("\n   �� SUCCESS! 100%% Accuracy Match with Python! ��\n");
        end else begin
            $display("\n   [FAIL] There were errors.\n");
        end
        $display("------------------------------------------------");
        $finish;
    end

endmodule