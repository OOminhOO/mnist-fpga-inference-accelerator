`timescale 1ns/1ps

module simple_score_overlay #(
    parameter H_VISIBLE = 640,
    parameter V_VISIBLE = 480
)(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [9:0]  x,
    input  wire [9:0]  y,
    input  wire [3:0]  number, // 0~9 (CNN ���)
    output reg         draw_on // 1�̸� ���� �ȼ���
);

    // ----------------------------------------------------
    // ����: ��ġ �� ũ��
    // ----------------------------------------------------
    localparam START_X = 32;  // ȭ�� �������� ������ �Ÿ�
    localparam START_Y = 32;  // ȭ�� ��ܿ��� ������ �Ÿ�
    localparam SCALE   = 4;   // ��Ʈ ũ�� Ȯ�� ���� (�⺻ 8x16 -> 32x64)
    
    // �⺻ ��Ʈ ũ�� (8x16)
    wire [3:0] font_col = (x - START_X) / SCALE; // 0..7
    wire [3:0] font_row = (y - START_Y) / SCALE; // 0..15

    // ���� ��ǥ�� ��Ʈ �ڽ� �ȿ� �ִ��� Ȯ��
    wire in_rect = (x >= START_X) && (x < START_X + 8*SCALE) &&
                   (y >= START_Y) && (y < START_Y + 16*SCALE);

    // ----------------------------------------------------
    // ��Ʈ ������ (0~9) - 8x16 ��Ʈ��
    // ----------------------------------------------------
    reg [7:0] font_data;
    
    always @(*) begin
        case ({number, font_row}) // {����, ��}
            // Number 0
            {4'd0, 4'd0 }: font_data = 8'h00; {4'd0, 4'd1 }: font_data = 8'h3C; {4'd0, 4'd2 }: font_data = 8'h42; {4'd0, 4'd3 }: font_data = 8'h42;
            {4'd0, 4'd4 }: font_data = 8'h42; {4'd0, 4'd5 }: font_data = 8'h42; {4'd0, 4'd6 }: font_data = 8'h42; {4'd0, 4'd7 }: font_data = 8'h42;
            {4'd0, 4'd8 }: font_data = 8'h42; {4'd0, 4'd9 }: font_data = 8'h42; {4'd0, 4'd10}: font_data = 8'h42; {4'd0, 4'd11}: font_data = 8'h42;
            {4'd0, 4'd12}: font_data = 8'h42; {4'd0, 4'd13}: font_data = 8'h42; {4'd0, 4'd14}: font_data = 8'h3C; {4'd0, 4'd15}: font_data = 8'h00;
            
            // Number 1
            {4'd1, 4'd0 }: font_data = 8'h00; {4'd1, 4'd1 }: font_data = 8'h08; {4'd1, 4'd2 }: font_data = 8'h18; {4'd1, 4'd3 }: font_data = 8'h28;
            {4'd1, 4'd4 }: font_data = 8'h08; {4'd1, 4'd5 }: font_data = 8'h08; {4'd1, 4'd6 }: font_data = 8'h08; {4'd1, 4'd7 }: font_data = 8'h08;
            {4'd1, 4'd8 }: font_data = 8'h08; {4'd1, 4'd9 }: font_data = 8'h08; {4'd1, 4'd10}: font_data = 8'h08; {4'd1, 4'd11}: font_data = 8'h08;
            {4'd1, 4'd12}: font_data = 8'h08; {4'd1, 4'd13}: font_data = 8'h08; {4'd1, 4'd14}: font_data = 8'h3E; {4'd0, 4'd15}: font_data = 8'h00;

            // Number 2
            {4'd2, 4'd0 }: font_data = 8'h00; {4'd2, 4'd1 }: font_data = 8'h3C; {4'd2, 4'd2 }: font_data = 8'h42; {4'd2, 4'd3 }: font_data = 8'h42;
            {4'd2, 4'd4 }: font_data = 8'h02; {4'd2, 4'd5 }: font_data = 8'h02; {4'd2, 4'd6 }: font_data = 8'h04; {4'd2, 4'd7 }: font_data = 8'h08;
            {4'd2, 4'd8 }: font_data = 8'h10; {4'd2, 4'd9 }: font_data = 8'h20; {4'd2, 4'd10}: font_data = 8'h40; {4'd2, 4'd11}: font_data = 8'h80;
            {4'd2, 4'd12}: font_data = 8'h80; {4'd2, 4'd13}: font_data = 8'h80; {4'd2, 4'd14}: font_data = 8'hFE; {4'd2, 4'd15}: font_data = 8'h00;

            // Number 3
            {4'd3, 4'd0 }: font_data = 8'h00; {4'd3, 4'd1 }: font_data = 8'h3C; {4'd3, 4'd2 }: font_data = 8'h42; {4'd3, 4'd3 }: font_data = 8'h42;
            {4'd3, 4'd4 }: font_data = 8'h02; {4'd3, 4'd5 }: font_data = 8'h02; {4'd3, 4'd6 }: font_data = 8'h1C; {4'd3, 4'd7 }: font_data = 8'h02;
            {4'd3, 4'd8 }: font_data = 8'h02; {4'd3, 4'd9 }: font_data = 8'h02; {4'd3, 4'd10}: font_data = 8'h02; {4'd3, 4'd11}: font_data = 8'h02;
            {4'd3, 4'd12}: font_data = 8'h42; {4'd3, 4'd13}: font_data = 8'h42; {4'd3, 4'd14}: font_data = 8'h3C; {4'd3, 4'd15}: font_data = 8'h00;

            // Number 4
            {4'd4, 4'd0 }: font_data = 8'h00; {4'd4, 4'd1 }: font_data = 8'h04; {4'd4, 4'd2 }: font_data = 8'h0C; {4'd4, 4'd3 }: font_data = 8'h14;
            {4'd4, 4'd4 }: font_data = 8'h24; {4'd4, 4'd5 }: font_data = 8'h44; {4'd4, 4'd6 }: font_data = 8'h44; {4'd4, 4'd7 }: font_data = 8'h84;
            {4'd4, 4'd8 }: font_data = 8'hFE; {4'd4, 4'd9 }: font_data = 8'h04; {4'd4, 4'd10}: font_data = 8'h04; {4'd4, 4'd11}: font_data = 8'h04;
            {4'd4, 4'd12}: font_data = 8'h04; {4'd4, 4'd13}: font_data = 8'h04; {4'd4, 4'd14}: font_data = 8'h04; {4'd4, 4'd15}: font_data = 8'h00;

            // Number 5
            {4'd5, 4'd0 }: font_data = 8'h00; {4'd5, 4'd1 }: font_data = 8'hFE; {4'd5, 4'd2 }: font_data = 8'h80; {4'd5, 4'd3 }: font_data = 8'h80;
            {4'd5, 4'd4 }: font_data = 8'h80; {4'd5, 4'd5 }: font_data = 8'hFC; {4'd5, 4'd6 }: font_data = 8'h02; {4'd5, 4'd7 }: font_data = 8'h02;
            {4'd5, 4'd8 }: font_data = 8'h02; {4'd5, 4'd9 }: font_data = 8'h02; {4'd5, 4'd10}: font_data = 8'h02; {4'd5, 4'd11}: font_data = 8'h02;
            {4'd5, 4'd12}: font_data = 8'h82; {4'd5, 4'd13}: font_data = 8'h42; {4'd5, 4'd14}: font_data = 8'h3C; {4'd5, 4'd15}: font_data = 8'h00;

            // Number 6
            {4'd6, 4'd0 }: font_data = 8'h00; {4'd6, 4'd1 }: font_data = 8'h3C; {4'd6, 4'd2 }: font_data = 8'h42; {4'd6, 4'd3 }: font_data = 8'h80;
            {4'd6, 4'd4 }: font_data = 8'h80; {4'd6, 4'd5 }: font_data = 8'h80; {4'd6, 4'd6 }: font_data = 8'hBC; {4'd6, 4'd7 }: font_data = 8'hC2;
            {4'd6, 4'd8 }: font_data = 8'h82; {4'd6, 4'd9 }: font_data = 8'h82; {4'd6, 4'd10}: font_data = 8'h82; {4'd6, 4'd11}: font_data = 8'h82;
            {4'd6, 4'd12}: font_data = 8'h42; {4'd6, 4'd13}: font_data = 8'h42; {4'd6, 4'd14}: font_data = 8'h3C; {4'd6, 4'd15}: font_data = 8'h00;

            // Number 7
            {4'd7, 4'd0 }: font_data = 8'h00; {4'd7, 4'd1 }: font_data = 8'hFE; {4'd7, 4'd2 }: font_data = 8'h02; {4'd7, 4'd3 }: font_data = 8'h04;
            {4'd7, 4'd4 }: font_data = 8'h04; {4'd7, 4'd5 }: font_data = 8'h08; {4'd7, 4'd6 }: font_data = 8'h08; {4'd7, 4'd7 }: font_data = 8'h10;
            {4'd7, 4'd8 }: font_data = 8'h10; {4'd7, 4'd9 }: font_data = 8'h20; {4'd7, 4'd10}: font_data = 8'h20; {4'd7, 4'd11}: font_data = 8'h20;
            {4'd7, 4'd12}: font_data = 8'h20; {4'd7, 4'd13}: font_data = 8'h20; {4'd7, 4'd14}: font_data = 8'h20; {4'd7, 4'd15}: font_data = 8'h00;

            // Number 8
            {4'd8, 4'd0 }: font_data = 8'h00; {4'd8, 4'd1 }: font_data = 8'h3C; {4'd8, 4'd2 }: font_data = 8'h42; {4'd8, 4'd3 }: font_data = 8'h42;
            {4'd8, 4'd4 }: font_data = 8'h42; {4'd8, 4'd5 }: font_data = 8'h42; {4'd8, 4'd6 }: font_data = 8'h3C; {4'd8, 4'd7 }: font_data = 8'h42;
            {4'd8, 4'd8 }: font_data = 8'h42; {4'd8, 4'd9 }: font_data = 8'h42; {4'd8, 4'd10}: font_data = 8'h42; {4'd8, 4'd11}: font_data = 8'h42;
            {4'd8, 4'd12}: font_data = 8'h42; {4'd8, 4'd13}: font_data = 8'h42; {4'd8, 4'd14}: font_data = 8'h3C; {4'd8, 4'd15}: font_data = 8'h00;

            // Number 9
            {4'd9, 4'd0 }: font_data = 8'h00; {4'd9, 4'd1 }: font_data = 8'h3C; {4'd9, 4'd2 }: font_data = 8'h42; {4'd9, 4'd3 }: font_data = 8'h42;
            {4'd9, 4'd4 }: font_data = 8'h42; {4'd9, 4'd5 }: font_data = 8'h42; {4'd9, 4'd6 }: font_data = 8'h46; {4'd9, 4'd7 }: font_data = 8'h3A;
            {4'd9, 4'd8 }: font_data = 8'h02; {4'd9, 4'd9 }: font_data = 8'h02; {4'd9, 4'd10}: font_data = 8'h02; {4'd9, 4'd11}: font_data = 8'h02;
            {4'd9, 4'd12}: font_data = 8'h42; {4'd9, 4'd13}: font_data = 8'h42; {4'd9, 4'd14}: font_data = 8'h3C; {4'd9, 4'd15}: font_data = 8'h00;
            
            default:      font_data = 8'h00;
        endcase
    end

    always @(posedge clk) begin
        if (in_rect) begin
            // 8��Ʈ ������ �� ���� x�� �ش��ϴ� ��Ʈ�� 1���� Ȯ�� (MSB first)
            draw_on <= font_data[7 - font_col]; 
        end else begin
            draw_on <= 1'b0;
        end
    end

endmodule