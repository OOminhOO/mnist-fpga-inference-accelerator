`timescale 1ns / 1ps

(* use_dsp = "no" *)
module fully_connected (
    input  wire               clk,
    input  wire               rst_n,
    
    input  wire               in_valid,
    input  wire [7:0]         in_1, // Ch0
    input  wire [7:0]         in_2, // Ch1
    input  wire [7:0]         in_3, // Ch2

    output reg                out_valid,
    output reg  [3:0]         out_cls,
    output reg  signed [31:0] out_logit,
    output reg                out_last
);

    // 1. �޸� �ε�
    reg signed [7:0]  w_mem [0:479];
    reg signed [31:0] b_mem [0:9];

    // �� ������ �κ�: ���� ��� ���
    initial begin
        $readmemh("Wd.txt", w_mem); 
        $readmemh("bd.txt", b_mem);
    end

    // 2. ���� ��ȣ �� ���������� ��������
    reg [4:0]  cnt_in;
    reg [3:0]  cnt_out;
    reg        calc_busy;
    reg        out_busy;

    // ���������� �������� ���� (Stage 0 -> Stage 1 -> Stage 2)
    reg        valid_st0;      // ����ġ �б� ��ȿ
    reg [4:0]  cnt_in_st0;     
    
    reg        valid_st1;      // ���� ��ȿ
    reg [4:0]  cnt_in_st1;

    // �Է� ������ ������ (����ġ �д� ���� ��ٷ��� ��)
    reg [7:0]  in_1_d, in_2_d, in_3_d;

    // ������
    reg signed [31:0] acc [0:9]; 

    // 3. ���������� ���� (10�� ����)
    genvar i;
    generate
        for (i = 0; i < 10; i = i + 1) begin : PE_ARRAY
            
            // [Stage 0] ����ġ �б� (Registering)
            reg signed [7:0] w1, w2, w3;
            
            always @(posedge clk) begin
                // cnt_in�� ���� �̸� �о��
                w1 <= w_mem[((cnt_in * 3) + 0) * 10 + i];
                w2 <= w_mem[((cnt_in * 3) + 1) * 10 + i];
                w3 <= w_mem[((cnt_in * 3) + 2) * 10 + i];
            end

            // [Stage 1] ���� (Multiplier)
            // w1, w2, w3�� �̹� 1Ŭ�� ���� cnt_in�� �ش��ϴ� ����.
            // ���� �Է� ������(in_1)�� 1Ŭ�� ������ ��(in_1_d)�� ��� ¦�� ����.
            reg signed [15:0] m1, m2, m3;

            always @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    m1 <= 0; m2 <= 0; m3 <= 0;
                end else if (valid_st0) begin
                    m1 <= $signed({1'b0, in_1_d}) * w1;
                    m2 <= $signed({1'b0, in_2_d}) * w2;
                    m3 <= $signed({1'b0, in_3_d}) * w3;
                end
            end

            // [Stage 2] ���� (Accumulate)
            // 16��Ʈ ���� ��� 3���� 32��Ʈ ��ȣ Ȯ��(Sign Extension) �� ����
            wire signed [31:0] sum_m;
            assign sum_m = {{16{m1[15]}}, m1} + {{16{m2[15]}}, m2} + {{16{m3[15]}}, m3};

            always @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    acc[i] <= 0;
                end else if (valid_st1) begin
                    if (cnt_in_st1 == 0) begin
                        // ù ��° ��: Bias + ���� ��
                        acc[i] <= b_mem[i] + sum_m;
                    end else begin
                        // �� ��: ���� Acc + ���� ��
                        acc[i] <= acc[i] + sum_m;
                    end
                end
            end
        end
    endgenerate

    // 4. ���� ����
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt_in <= 0; 
            valid_st0 <= 0; cnt_in_st0 <= 0;
            valid_st1 <= 0; cnt_in_st1 <= 0;
            
            cnt_out <= 0; calc_busy <= 0; out_busy <= 0;
            out_valid <= 0; out_last <= 0; out_cls <= 0; out_logit <= 0;
            
            in_1_d <= 0; in_2_d <= 0; in_3_d <= 0;
        end else begin
            // [�Է� ����������]
            if (in_valid) begin
                calc_busy  <= 1;
                
                // Stage 0���� �ѱ�� ��ȣ
                valid_st0  <= 1;
                cnt_in_st0 <= cnt_in;
                
                // �Է� �����͵� 1Ŭ�� ������ (����ġ �д� �ð��� ����ȭ)
                in_1_d <= in_1;
                in_2_d <= in_2;
                in_3_d <= in_3;

                if (cnt_in == 15) begin
                    cnt_in <= 0;
                    calc_busy <= 0;
                end else begin
                    cnt_in <= cnt_in + 1;
                end
            end else begin
                valid_st0 <= 0;
            end

            // [Stage 0 -> Stage 1]
            valid_st1  <= valid_st0;
            cnt_in_st1 <= cnt_in_st0;

            // [��� Ÿ�̹�]
            // cnt_in_st1�� 15�̰�, valid_st1�� 1�̸� -> Stage 2���� ������ ���� �Ϸ��
            if (valid_st1 && (cnt_in_st1 == 15)) begin
                out_busy <= 1;
                cnt_out  <= 0;
            end

            // [��� ���]
            if (out_busy) begin
                out_valid <= 1;
                out_cls   <= cnt_out;
                out_logit <= acc[cnt_out]; 

                if (cnt_out == 9) begin
                    out_last <= 1;
                    out_busy <= 0;
                    cnt_out  <= 0;
                end else begin
                    out_last <= 0;
                    cnt_out  <= cnt_out + 1;
                end
            end else begin
                out_valid <= 0;
                out_last  <= 0;
            end
        end
    end

endmodule