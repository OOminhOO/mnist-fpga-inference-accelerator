`timescale 1ns / 1ps

module comparator (
    input  wire               clk,
    input  wire               rst_n,
    input  wire               in_valid,
    // in_sof ���� (in_cls == 0 ���� �Ǵ�)
    input  wire [3:0]         in_cls,
    input  wire signed [31:0] in_logit,
    input  wire               in_last,

    output reg  [3:0]         decision,
    output reg                out_valid
);
    reg signed [31:0] best_logit;
    reg [3:0]         best_cls;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            best_logit <= -32'sd2147483648; // �ּҰ� (Signed 32bit Min)
            best_cls   <= 4'd0;
            decision   <= 4'd0;
            out_valid  <= 1'b0;
        end else begin
            out_valid <= 1'b0; // ��ҿ� 0 (Pulse)

            if (in_valid) begin
                // 1. ù ��° Ŭ����(0��)�� ������ ������ �ʱ�ȭ
                if (in_cls == 4'd0) begin
                    best_logit <= in_logit;
                    best_cls   <= in_cls;
                end 
                // 2. �� �� (1~9��): ���� ���� �� ũ�� ����
                else begin
                    if (in_logit > best_logit) begin
                        best_logit <= in_logit;
                        best_cls   <= in_cls;
                    end
                end

                // 3. ������ Ŭ����(9��)�� �� ���� ���� (Ÿ�̹� ���� ����)
                if (in_last) begin
                    out_valid <= 1'b1;
                    
                    // �� �߿�: 9���� ���� 1��� ũ�� 9���� ���, �ƴϸ� ���� 1�� ���
                    // (best_logit�� ���� ������Ʈ �Ǳ� �� ���� ������ �����Ƿ� ���⼭ ���ؾ� ��)
                    if (in_cls == 4'd0) begin
                        // Ȥ�ö� Ŭ������ 1������ ��� (����ڵ�)
                        decision <= in_cls;
                    end 
                    else if (in_logit > best_logit) begin
                        decision <= in_cls; // ��� ���� 9���� ������!
                    end else begin
                        decision <= best_cls; // ���� 1�� ����
                    end
                end
            end
        end
    end
endmodule